*A BUS interconnect circuit with 10 bus line 8 segment.

Rin1 0 TDn1a1 10
Rin2 0 TDn2a1 10
Rin3 0 TDn3a1 10
Rin4 0 TDn4a1 10
Rin5 0 TDn5a1 10
Rin6 0 TDn6a1 10
Rin7 0 TDn7a1 10
Rin8 0 TDn8a1 10
*Iin1 TDn1a1 0 AC 1
Iin1 TDn1a1 0 PULSE(0 1 0.05ns 0.05ns 0.05ns 0.30ns 0.50ns)

Rgndg TDnga1 0 1
Rvndg TDnva1 0 1
RRR TDnga9 TDnva9 1
Cout1 TDn1a9 TDnga9 0.1p
Cout2 TDn2a9 TDnga9 0.1p
Cout3 TDn3a9 TDnga9 0.1p
Cout4 TDn4a9 TDnga9 0.1p
Cout5 TDn5a9 TDnga9 0.1p
Cout6 TDn6a9 TDnga9 0.1p
Cout7 TDn7a9 TDnga9 0.1p
Cout8 TDn8a9 TDnga9 0.1p

X1 TDnga1 TDnga9 TDn1a1 TDn1a9 TDn2a1 TDn2a9 TDn3a1 TDn3a9 TDn4a1 TDn4a9 TDn5a1 TDn5a9 TDn6a1 TDn6a9 TDn7a1 TDn7a9 TDn8a1 TDn8a9 TDnva1 TDnva9 intercon
.SUBCKT intercon TDnga1 TDnga17 TDn1a1 TDn1a17 TDn2a1 TDn2a17 TDn3a1 TDn3a17 TDn4a1 TDn4a17 TDn5a1 TDn5a17 TDn6a1 TDn6a17 TDn7a1 TDn7a17 TDn8a1 TDn8a17 TDnva1 TDnva17

Rnga1 TDnga1 TDnga2 2.603750
Rnga2 TDnga3 TDnga4 2.603750
Rnga3 TDnga5 TDnga6 2.603750
Rnga4 TDnga7 TDnga8 2.603750
Rnga5 TDnga9 TDnga10 2.603750
Rnga6 TDnga11 TDnga12 2.603750
Rnga7 TDnga13 TDnga14 2.603750
Rnga8 TDnga15 TDnga16 2.603750
Rn1a1 TDn1a1 TDn1a2 2.604380
Rn1a2 TDn1a3 TDn1a4 2.604380
Rn1a3 TDn1a5 TDn1a6 2.604380
Rn1a4 TDn1a7 TDn1a8 2.604380
Rn1a5 TDn1a9 TDn1a10 2.604380
Rn1a6 TDn1a11 TDn1a12 2.604380
Rn1a7 TDn1a13 TDn1a14 2.604380
Rn1a8 TDn1a15 TDn1a16 2.604380
Rn2a1 TDn2a1 TDn2a2 2.604380
Rn2a2 TDn2a3 TDn2a4 2.604380
Rn2a3 TDn2a5 TDn2a6 2.604380
Rn2a4 TDn2a7 TDn2a8 2.604380
Rn2a5 TDn2a9 TDn2a10 2.604380
Rn2a6 TDn2a11 TDn2a12 2.604380
Rn2a7 TDn2a13 TDn2a14 2.604380
Rn2a8 TDn2a15 TDn2a16 2.604380
Rn3a1 TDn3a1 TDn3a2 2.604380
Rn3a2 TDn3a3 TDn3a4 2.604380
Rn3a3 TDn3a5 TDn3a6 2.604380
Rn3a4 TDn3a7 TDn3a8 2.604380
Rn3a5 TDn3a9 TDn3a10 2.604380
Rn3a6 TDn3a11 TDn3a12 2.604380
Rn3a7 TDn3a13 TDn3a14 2.604380
Rn3a8 TDn3a15 TDn3a16 2.604380
Rn4a1 TDn4a1 TDn4a2 2.604380
Rn4a2 TDn4a3 TDn4a4 2.604380
Rn4a3 TDn4a5 TDn4a6 2.604380
Rn4a4 TDn4a7 TDn4a8 2.604380
Rn4a5 TDn4a9 TDn4a10 2.604380
Rn4a6 TDn4a11 TDn4a12 2.604380
Rn4a7 TDn4a13 TDn4a14 2.604380
Rn4a8 TDn4a15 TDn4a16 2.604380
Rn5a1 TDn5a1 TDn5a2 2.604380
Rn5a2 TDn5a3 TDn5a4 2.604380
Rn5a3 TDn5a5 TDn5a6 2.604380
Rn5a4 TDn5a7 TDn5a8 2.604380
Rn5a5 TDn5a9 TDn5a10 2.604380
Rn5a6 TDn5a11 TDn5a12 2.604380
Rn5a7 TDn5a13 TDn5a14 2.604380
Rn5a8 TDn5a15 TDn5a16 2.604380
Rn6a1 TDn6a1 TDn6a2 2.604380
Rn6a2 TDn6a3 TDn6a4 2.604380
Rn6a3 TDn6a5 TDn6a6 2.604380
Rn6a4 TDn6a7 TDn6a8 2.604380
Rn6a5 TDn6a9 TDn6a10 2.604380
Rn6a6 TDn6a11 TDn6a12 2.604380
Rn6a7 TDn6a13 TDn6a14 2.604380
Rn6a8 TDn6a15 TDn6a16 2.604380
Rn7a1 TDn7a1 TDn7a2 2.604380
Rn7a2 TDn7a3 TDn7a4 2.604380
Rn7a3 TDn7a5 TDn7a6 2.604380
Rn7a4 TDn7a7 TDn7a8 2.604380
Rn7a5 TDn7a9 TDn7a10 2.604380
Rn7a6 TDn7a11 TDn7a12 2.604380
Rn7a7 TDn7a13 TDn7a14 2.604380
Rn7a8 TDn7a15 TDn7a16 2.604380
Rn8a1 TDn8a1 TDn8a2 2.604380
Rn8a2 TDn8a3 TDn8a4 2.604380
Rn8a3 TDn8a5 TDn8a6 2.604380
Rn8a4 TDn8a7 TDn8a8 2.604380
Rn8a5 TDn8a9 TDn8a10 2.604380
Rn8a6 TDn8a11 TDn8a12 2.604380
Rn8a7 TDn8a13 TDn8a14 2.604380
Rn8a8 TDn8a15 TDn8a16 2.604380
Rnva1 TDnva1 TDnva2 2.603750
Rnva2 TDnva3 TDnva4 2.603750
Rnva3 TDnva5 TDnva6 2.603750
Rnva4 TDnva7 TDnva8 2.603750
Rnva5 TDnva9 TDnva10 2.603750
Rnva6 TDnva11 TDnva12 2.603750
Rnva7 TDnva13 TDnva14 2.603750
Rnva8 TDnva15 TDnva16 2.603750
Lnga1 TDnga2 TDnga3 8.243750e-010
Lnga2 TDnga4 TDnga5 8.243750e-010
Lnga3 TDnga6 TDnga7 8.243750e-010
Lnga4 TDnga8 TDnga9 8.243750e-010
Lnga5 TDnga10 TDnga11 8.243750e-010
Lnga6 TDnga12 TDnga13 8.243750e-010
Lnga7 TDnga14 TDnga15 8.243750e-010
Lnga8 TDnga16 TDnga17 8.243750e-010
Ln1a1 TDn1a2 TDn1a3 8.243750e-010
Ln1a2 TDn1a4 TDn1a5 8.243750e-010
Ln1a3 TDn1a6 TDn1a7 8.243750e-010
Ln1a4 TDn1a8 TDn1a9 8.243750e-010
Ln1a5 TDn1a10 TDn1a11 8.243750e-010
Ln1a6 TDn1a12 TDn1a13 8.243750e-010
Ln1a7 TDn1a14 TDn1a15 8.243750e-010
Ln1a8 TDn1a16 TDn1a17 8.243750e-010
Ln2a1 TDn2a2 TDn2a3 8.243750e-010
Ln2a2 TDn2a4 TDn2a5 8.243750e-010
Ln2a3 TDn2a6 TDn2a7 8.243750e-010
Ln2a4 TDn2a8 TDn2a9 8.243750e-010
Ln2a5 TDn2a10 TDn2a11 8.243750e-010
Ln2a6 TDn2a12 TDn2a13 8.243750e-010
Ln2a7 TDn2a14 TDn2a15 8.243750e-010
Ln2a8 TDn2a16 TDn2a17 8.243750e-010
Ln3a1 TDn3a2 TDn3a3 8.243750e-010
Ln3a2 TDn3a4 TDn3a5 8.243750e-010
Ln3a3 TDn3a6 TDn3a7 8.243750e-010
Ln3a4 TDn3a8 TDn3a9 8.243750e-010
Ln3a5 TDn3a10 TDn3a11 8.243750e-010
Ln3a6 TDn3a12 TDn3a13 8.243750e-010
Ln3a7 TDn3a14 TDn3a15 8.243750e-010
Ln3a8 TDn3a16 TDn3a17 8.243750e-010
Ln4a1 TDn4a2 TDn4a3 8.243750e-010
Ln4a2 TDn4a4 TDn4a5 8.243750e-010
Ln4a3 TDn4a6 TDn4a7 8.243750e-010
Ln4a4 TDn4a8 TDn4a9 8.243750e-010
Ln4a5 TDn4a10 TDn4a11 8.243750e-010
Ln4a6 TDn4a12 TDn4a13 8.243750e-010
Ln4a7 TDn4a14 TDn4a15 8.243750e-010
Ln4a8 TDn4a16 TDn4a17 8.243750e-010
Ln5a1 TDn5a2 TDn5a3 8.243750e-010
Ln5a2 TDn5a4 TDn5a5 8.243750e-010
Ln5a3 TDn5a6 TDn5a7 8.243750e-010
Ln5a4 TDn5a8 TDn5a9 8.243750e-010
Ln5a5 TDn5a10 TDn5a11 8.243750e-010
Ln5a6 TDn5a12 TDn5a13 8.243750e-010
Ln5a7 TDn5a14 TDn5a15 8.243750e-010
Ln5a8 TDn5a16 TDn5a17 8.243750e-010
Ln6a1 TDn6a2 TDn6a3 8.243750e-010
Ln6a2 TDn6a4 TDn6a5 8.243750e-010
Ln6a3 TDn6a6 TDn6a7 8.243750e-010
Ln6a4 TDn6a8 TDn6a9 8.243750e-010
Ln6a5 TDn6a10 TDn6a11 8.243750e-010
Ln6a6 TDn6a12 TDn6a13 8.243750e-010
Ln6a7 TDn6a14 TDn6a15 8.243750e-010
Ln6a8 TDn6a16 TDn6a17 8.243750e-010
Ln7a1 TDn7a2 TDn7a3 8.243750e-010
Ln7a2 TDn7a4 TDn7a5 8.243750e-010
Ln7a3 TDn7a6 TDn7a7 8.243750e-010
Ln7a4 TDn7a8 TDn7a9 8.243750e-010
Ln7a5 TDn7a10 TDn7a11 8.243750e-010
Ln7a6 TDn7a12 TDn7a13 8.243750e-010
Ln7a7 TDn7a14 TDn7a15 8.243750e-010
Ln7a8 TDn7a16 TDn7a17 8.243750e-010
Ln8a1 TDn8a2 TDn8a3 8.243750e-010
Ln8a2 TDn8a4 TDn8a5 8.243750e-010
Ln8a3 TDn8a6 TDn8a7 8.243750e-010
Ln8a4 TDn8a8 TDn8a9 8.243750e-010
Ln8a5 TDn8a10 TDn8a11 8.243750e-010
Ln8a6 TDn8a12 TDn8a13 8.243750e-010
Ln8a7 TDn8a14 TDn8a15 8.243750e-010
Ln8a8 TDn8a16 TDn8a17 8.243750e-010
Lnva1 TDnva2 TDnva3 8.243750e-010
Lnva2 TDnva4 TDnva5 8.243750e-010
Lnva3 TDnva6 TDnva7 8.243750e-010
Lnva4 TDnva8 TDnva9 8.243750e-010
Lnva5 TDnva10 TDnva11 8.243750e-010
Lnva6 TDnva12 TDnva13 8.243750e-010
Lnva7 TDnva14 TDnva15 8.243750e-010
Lnva8 TDnva16 TDnva17 8.243750e-010
Kngan1a1 Lnga1 Ln1a1 0.805155
Kngan1a2 Lnga2 Ln1a2 0.805155
Kngan1a3 Lnga3 Ln1a3 0.805155
Kngan1a4 Lnga4 Ln1a4 0.805155
Kngan1a5 Lnga5 Ln1a5 0.805155
Kngan1a6 Lnga6 Ln1a6 0.805155
Kngan1a7 Lnga7 Ln1a7 0.805155
Kngan1a8 Lnga8 Ln1a8 0.805155
Kngan2a1 Lnga1 Ln2a1 0.723730
Kngan2a2 Lnga2 Ln2a2 0.723730
Kngan2a3 Lnga3 Ln2a3 0.723730
Kngan2a4 Lnga4 Ln2a4 0.723730
Kngan2a5 Lnga5 Ln2a5 0.723730
Kngan2a6 Lnga6 Ln2a6 0.723730
Kngan2a7 Lnga7 Ln2a7 0.723730
Kngan2a8 Lnga8 Ln2a8 0.723730
Kngan3a1 Lnga1 Ln3a1 0.675208
Kngan3a2 Lnga2 Ln3a2 0.675208
Kngan3a3 Lnga3 Ln3a3 0.675208
Kngan3a4 Lnga4 Ln3a4 0.675208
Kngan3a5 Lnga5 Ln3a5 0.675208
Kngan3a6 Lnga6 Ln3a6 0.675208
Kngan3a7 Lnga7 Ln3a7 0.675208
Kngan3a8 Lnga8 Ln3a8 0.675208
Kngan4a1 Lnga1 Ln4a1 0.640637
Kngan4a2 Lnga2 Ln4a2 0.640637
Kngan4a3 Lnga3 Ln4a3 0.640637
Kngan4a4 Lnga4 Ln4a4 0.640637
Kngan4a5 Lnga5 Ln4a5 0.640637
Kngan4a6 Lnga6 Ln4a6 0.640637
Kngan4a7 Lnga7 Ln4a7 0.640637
Kngan4a8 Lnga8 Ln4a8 0.640637
Kngan5a1 Lnga1 Ln5a1 0.613723
Kngan5a2 Lnga2 Ln5a2 0.613723
Kngan5a3 Lnga3 Ln5a3 0.613723
Kngan5a4 Lnga4 Ln5a4 0.613723
Kngan5a5 Lnga5 Ln5a5 0.613723
Kngan5a6 Lnga6 Ln5a6 0.613723
Kngan5a7 Lnga7 Ln5a7 0.613723
Kngan5a8 Lnga8 Ln5a8 0.613723
Kngan6a1 Lnga1 Ln6a1 0.591812
Kngan6a2 Lnga2 Ln6a2 0.591812
Kngan6a3 Lnga3 Ln6a3 0.591812
Kngan6a4 Lnga4 Ln6a4 0.591812
Kngan6a5 Lnga5 Ln6a5 0.591812
Kngan6a6 Lnga6 Ln6a6 0.591812
Kngan6a7 Lnga7 Ln6a7 0.591812
Kngan6a8 Lnga8 Ln6a8 0.591812
Kngan7a1 Lnga1 Ln7a1 0.573237
Kngan7a2 Lnga2 Ln7a2 0.573237
Kngan7a3 Lnga3 Ln7a3 0.573237
Kngan7a4 Lnga4 Ln7a4 0.573237
Kngan7a5 Lnga5 Ln7a5 0.573237
Kngan7a6 Lnga6 Ln7a6 0.573237
Kngan7a7 Lnga7 Ln7a7 0.573237
Kngan7a8 Lnga8 Ln7a8 0.573237
Kngan8a1 Lnga1 Ln8a1 0.557165
Kngan8a2 Lnga2 Ln8a2 0.557165
Kngan8a3 Lnga3 Ln8a3 0.557165
Kngan8a4 Lnga4 Ln8a4 0.557165
Kngan8a5 Lnga5 Ln8a5 0.557165
Kngan8a6 Lnga6 Ln8a6 0.557165
Kngan8a7 Lnga7 Ln8a7 0.557165
Kngan8a8 Lnga8 Ln8a8 0.557165
Knganva1 Lnga1 Lnva1 0.542987
Knganva2 Lnga2 Lnva2 0.542987
Knganva3 Lnga3 Lnva3 0.542987
Knganva4 Lnga4 Lnva4 0.542987
Knganva5 Lnga5 Lnva5 0.542987
Knganva6 Lnga6 Lnva6 0.542987
Knganva7 Lnga7 Lnva7 0.542987
Knganva8 Lnga8 Lnva8 0.542987
Kn1an2a1 Ln1a1 Ln2a1 0.805155
Kn1an2a2 Ln1a2 Ln2a2 0.805155
Kn1an2a3 Ln1a3 Ln2a3 0.805155
Kn1an2a4 Ln1a4 Ln2a4 0.805155
Kn1an2a5 Ln1a5 Ln2a5 0.805155
Kn1an2a6 Ln1a6 Ln2a6 0.805155
Kn1an2a7 Ln1a7 Ln2a7 0.805155
Kn1an2a8 Ln1a8 Ln2a8 0.805155
Kn1an3a1 Ln1a1 Ln3a1 0.723730
Kn1an3a2 Ln1a2 Ln3a2 0.723730
Kn1an3a3 Ln1a3 Ln3a3 0.723730
Kn1an3a4 Ln1a4 Ln3a4 0.723730
Kn1an3a5 Ln1a5 Ln3a5 0.723730
Kn1an3a6 Ln1a6 Ln3a6 0.723730
Kn1an3a7 Ln1a7 Ln3a7 0.723730
Kn1an3a8 Ln1a8 Ln3a8 0.723730
Kn1an4a1 Ln1a1 Ln4a1 0.675208
Kn1an4a2 Ln1a2 Ln4a2 0.675208
Kn1an4a3 Ln1a3 Ln4a3 0.675208
Kn1an4a4 Ln1a4 Ln4a4 0.675208
Kn1an4a5 Ln1a5 Ln4a5 0.675208
Kn1an4a6 Ln1a6 Ln4a6 0.675208
Kn1an4a7 Ln1a7 Ln4a7 0.675208
Kn1an4a8 Ln1a8 Ln4a8 0.675208
Kn1an5a1 Ln1a1 Ln5a1 0.640637
Kn1an5a2 Ln1a2 Ln5a2 0.640637
Kn1an5a3 Ln1a3 Ln5a3 0.640637
Kn1an5a4 Ln1a4 Ln5a4 0.640637
Kn1an5a5 Ln1a5 Ln5a5 0.640637
Kn1an5a6 Ln1a6 Ln5a6 0.640637
Kn1an5a7 Ln1a7 Ln5a7 0.640637
Kn1an5a8 Ln1a8 Ln5a8 0.640637
Kn1an6a1 Ln1a1 Ln6a1 0.613723
Kn1an6a2 Ln1a2 Ln6a2 0.613723
Kn1an6a3 Ln1a3 Ln6a3 0.613723
Kn1an6a4 Ln1a4 Ln6a4 0.613723
Kn1an6a5 Ln1a5 Ln6a5 0.613723
Kn1an6a6 Ln1a6 Ln6a6 0.613723
Kn1an6a7 Ln1a7 Ln6a7 0.613723
Kn1an6a8 Ln1a8 Ln6a8 0.613723
Kn1an7a1 Ln1a1 Ln7a1 0.591812
Kn1an7a2 Ln1a2 Ln7a2 0.591812
Kn1an7a3 Ln1a3 Ln7a3 0.591812
Kn1an7a4 Ln1a4 Ln7a4 0.591812
Kn1an7a5 Ln1a5 Ln7a5 0.591812
Kn1an7a6 Ln1a6 Ln7a6 0.591812
Kn1an7a7 Ln1a7 Ln7a7 0.591812
Kn1an7a8 Ln1a8 Ln7a8 0.591812
Kn1an8a1 Ln1a1 Ln8a1 0.573237
Kn1an8a2 Ln1a2 Ln8a2 0.573237
Kn1an8a3 Ln1a3 Ln8a3 0.573237
Kn1an8a4 Ln1a4 Ln8a4 0.573237
Kn1an8a5 Ln1a5 Ln8a5 0.573237
Kn1an8a6 Ln1a6 Ln8a6 0.573237
Kn1an8a7 Ln1a7 Ln8a7 0.573237
Kn1an8a8 Ln1a8 Ln8a8 0.573237
Kn1anva1 Ln1a1 Lnva1 0.557165
Kn1anva2 Ln1a2 Lnva2 0.557165
Kn1anva3 Ln1a3 Lnva3 0.557165
Kn1anva4 Ln1a4 Lnva4 0.557165
Kn1anva5 Ln1a5 Lnva5 0.557165
Kn1anva6 Ln1a6 Lnva6 0.557165
Kn1anva7 Ln1a7 Lnva7 0.557165
Kn1anva8 Ln1a8 Lnva8 0.557165
Kn2an3a1 Ln2a1 Ln3a1 0.805155
Kn2an3a2 Ln2a2 Ln3a2 0.805155
Kn2an3a3 Ln2a3 Ln3a3 0.805155
Kn2an3a4 Ln2a4 Ln3a4 0.805155
Kn2an3a5 Ln2a5 Ln3a5 0.805155
Kn2an3a6 Ln2a6 Ln3a6 0.805155
Kn2an3a7 Ln2a7 Ln3a7 0.805155
Kn2an3a8 Ln2a8 Ln3a8 0.805155
Kn2an4a1 Ln2a1 Ln4a1 0.723730
Kn2an4a2 Ln2a2 Ln4a2 0.723730
Kn2an4a3 Ln2a3 Ln4a3 0.723730
Kn2an4a4 Ln2a4 Ln4a4 0.723730
Kn2an4a5 Ln2a5 Ln4a5 0.723730
Kn2an4a6 Ln2a6 Ln4a6 0.723730
Kn2an4a7 Ln2a7 Ln4a7 0.723730
Kn2an4a8 Ln2a8 Ln4a8 0.723730
Kn2an5a1 Ln2a1 Ln5a1 0.675208
Kn2an5a2 Ln2a2 Ln5a2 0.675208
Kn2an5a3 Ln2a3 Ln5a3 0.675208
Kn2an5a4 Ln2a4 Ln5a4 0.675208
Kn2an5a5 Ln2a5 Ln5a5 0.675208
Kn2an5a6 Ln2a6 Ln5a6 0.675208
Kn2an5a7 Ln2a7 Ln5a7 0.675208
Kn2an5a8 Ln2a8 Ln5a8 0.675208
Kn2an6a1 Ln2a1 Ln6a1 0.640637
Kn2an6a2 Ln2a2 Ln6a2 0.640637
Kn2an6a3 Ln2a3 Ln6a3 0.640637
Kn2an6a4 Ln2a4 Ln6a4 0.640637
Kn2an6a5 Ln2a5 Ln6a5 0.640637
Kn2an6a6 Ln2a6 Ln6a6 0.640637
Kn2an6a7 Ln2a7 Ln6a7 0.640637
Kn2an6a8 Ln2a8 Ln6a8 0.640637
Kn2an7a1 Ln2a1 Ln7a1 0.613723
Kn2an7a2 Ln2a2 Ln7a2 0.613723
Kn2an7a3 Ln2a3 Ln7a3 0.613723
Kn2an7a4 Ln2a4 Ln7a4 0.613723
Kn2an7a5 Ln2a5 Ln7a5 0.613723
Kn2an7a6 Ln2a6 Ln7a6 0.613723
Kn2an7a7 Ln2a7 Ln7a7 0.613723
Kn2an7a8 Ln2a8 Ln7a8 0.613723
Kn2an8a1 Ln2a1 Ln8a1 0.591812
Kn2an8a2 Ln2a2 Ln8a2 0.591812
Kn2an8a3 Ln2a3 Ln8a3 0.591812
Kn2an8a4 Ln2a4 Ln8a4 0.591812
Kn2an8a5 Ln2a5 Ln8a5 0.591812
Kn2an8a6 Ln2a6 Ln8a6 0.591812
Kn2an8a7 Ln2a7 Ln8a7 0.591812
Kn2an8a8 Ln2a8 Ln8a8 0.591812
Kn2anva1 Ln2a1 Lnva1 0.573237
Kn2anva2 Ln2a2 Lnva2 0.573237
Kn2anva3 Ln2a3 Lnva3 0.573237
Kn2anva4 Ln2a4 Lnva4 0.573237
Kn2anva5 Ln2a5 Lnva5 0.573237
Kn2anva6 Ln2a6 Lnva6 0.573237
Kn2anva7 Ln2a7 Lnva7 0.573237
Kn2anva8 Ln2a8 Lnva8 0.573237
Kn3an4a1 Ln3a1 Ln4a1 0.805155
Kn3an4a2 Ln3a2 Ln4a2 0.805155
Kn3an4a3 Ln3a3 Ln4a3 0.805155
Kn3an4a4 Ln3a4 Ln4a4 0.805155
Kn3an4a5 Ln3a5 Ln4a5 0.805155
Kn3an4a6 Ln3a6 Ln4a6 0.805155
Kn3an4a7 Ln3a7 Ln4a7 0.805155
Kn3an4a8 Ln3a8 Ln4a8 0.805155
Kn3an5a1 Ln3a1 Ln5a1 0.723730
Kn3an5a2 Ln3a2 Ln5a2 0.723730
Kn3an5a3 Ln3a3 Ln5a3 0.723730
Kn3an5a4 Ln3a4 Ln5a4 0.723730
Kn3an5a5 Ln3a5 Ln5a5 0.723730
Kn3an5a6 Ln3a6 Ln5a6 0.723730
Kn3an5a7 Ln3a7 Ln5a7 0.723730
Kn3an5a8 Ln3a8 Ln5a8 0.723730
Kn3an6a1 Ln3a1 Ln6a1 0.675208
Kn3an6a2 Ln3a2 Ln6a2 0.675208
Kn3an6a3 Ln3a3 Ln6a3 0.675208
Kn3an6a4 Ln3a4 Ln6a4 0.675208
Kn3an6a5 Ln3a5 Ln6a5 0.675208
Kn3an6a6 Ln3a6 Ln6a6 0.675208
Kn3an6a7 Ln3a7 Ln6a7 0.675208
Kn3an6a8 Ln3a8 Ln6a8 0.675208
Kn3an7a1 Ln3a1 Ln7a1 0.640637
Kn3an7a2 Ln3a2 Ln7a2 0.640637
Kn3an7a3 Ln3a3 Ln7a3 0.640637
Kn3an7a4 Ln3a4 Ln7a4 0.640637
Kn3an7a5 Ln3a5 Ln7a5 0.640637
Kn3an7a6 Ln3a6 Ln7a6 0.640637
Kn3an7a7 Ln3a7 Ln7a7 0.640637
Kn3an7a8 Ln3a8 Ln7a8 0.640637
Kn3an8a1 Ln3a1 Ln8a1 0.613723
Kn3an8a2 Ln3a2 Ln8a2 0.613723
Kn3an8a3 Ln3a3 Ln8a3 0.613723
Kn3an8a4 Ln3a4 Ln8a4 0.613723
Kn3an8a5 Ln3a5 Ln8a5 0.613723
Kn3an8a6 Ln3a6 Ln8a6 0.613723
Kn3an8a7 Ln3a7 Ln8a7 0.613723
Kn3an8a8 Ln3a8 Ln8a8 0.613723
Kn3anva1 Ln3a1 Lnva1 0.591812
Kn3anva2 Ln3a2 Lnva2 0.591812
Kn3anva3 Ln3a3 Lnva3 0.591812
Kn3anva4 Ln3a4 Lnva4 0.591812
Kn3anva5 Ln3a5 Lnva5 0.591812
Kn3anva6 Ln3a6 Lnva6 0.591812
Kn3anva7 Ln3a7 Lnva7 0.591812
Kn3anva8 Ln3a8 Lnva8 0.591812
Kn4an5a1 Ln4a1 Ln5a1 0.805155
Kn4an5a2 Ln4a2 Ln5a2 0.805155
Kn4an5a3 Ln4a3 Ln5a3 0.805155
Kn4an5a4 Ln4a4 Ln5a4 0.805155
Kn4an5a5 Ln4a5 Ln5a5 0.805155
Kn4an5a6 Ln4a6 Ln5a6 0.805155
Kn4an5a7 Ln4a7 Ln5a7 0.805155
Kn4an5a8 Ln4a8 Ln5a8 0.805155
Kn4an6a1 Ln4a1 Ln6a1 0.723730
Kn4an6a2 Ln4a2 Ln6a2 0.723730
Kn4an6a3 Ln4a3 Ln6a3 0.723730
Kn4an6a4 Ln4a4 Ln6a4 0.723730
Kn4an6a5 Ln4a5 Ln6a5 0.723730
Kn4an6a6 Ln4a6 Ln6a6 0.723730
Kn4an6a7 Ln4a7 Ln6a7 0.723730
Kn4an6a8 Ln4a8 Ln6a8 0.723730
Kn4an7a1 Ln4a1 Ln7a1 0.675208
Kn4an7a2 Ln4a2 Ln7a2 0.675208
Kn4an7a3 Ln4a3 Ln7a3 0.675208
Kn4an7a4 Ln4a4 Ln7a4 0.675208
Kn4an7a5 Ln4a5 Ln7a5 0.675208
Kn4an7a6 Ln4a6 Ln7a6 0.675208
Kn4an7a7 Ln4a7 Ln7a7 0.675208
Kn4an7a8 Ln4a8 Ln7a8 0.675208
Kn4an8a1 Ln4a1 Ln8a1 0.640637
Kn4an8a2 Ln4a2 Ln8a2 0.640637
Kn4an8a3 Ln4a3 Ln8a3 0.640637
Kn4an8a4 Ln4a4 Ln8a4 0.640637
Kn4an8a5 Ln4a5 Ln8a5 0.640637
Kn4an8a6 Ln4a6 Ln8a6 0.640637
Kn4an8a7 Ln4a7 Ln8a7 0.640637
Kn4an8a8 Ln4a8 Ln8a8 0.640637
Kn4anva1 Ln4a1 Lnva1 0.613723
Kn4anva2 Ln4a2 Lnva2 0.613723
Kn4anva3 Ln4a3 Lnva3 0.613723
Kn4anva4 Ln4a4 Lnva4 0.613723
Kn4anva5 Ln4a5 Lnva5 0.613723
Kn4anva6 Ln4a6 Lnva6 0.613723
Kn4anva7 Ln4a7 Lnva7 0.613723
Kn4anva8 Ln4a8 Lnva8 0.613723
Kn5an6a1 Ln5a1 Ln6a1 0.805155
Kn5an6a2 Ln5a2 Ln6a2 0.805155
Kn5an6a3 Ln5a3 Ln6a3 0.805155
Kn5an6a4 Ln5a4 Ln6a4 0.805155
Kn5an6a5 Ln5a5 Ln6a5 0.805155
Kn5an6a6 Ln5a6 Ln6a6 0.805155
Kn5an6a7 Ln5a7 Ln6a7 0.805155
Kn5an6a8 Ln5a8 Ln6a8 0.805155
Kn5an7a1 Ln5a1 Ln7a1 0.723730
Kn5an7a2 Ln5a2 Ln7a2 0.723730
Kn5an7a3 Ln5a3 Ln7a3 0.723730
Kn5an7a4 Ln5a4 Ln7a4 0.723730
Kn5an7a5 Ln5a5 Ln7a5 0.723730
Kn5an7a6 Ln5a6 Ln7a6 0.723730
Kn5an7a7 Ln5a7 Ln7a7 0.723730
Kn5an7a8 Ln5a8 Ln7a8 0.723730
Kn5an8a1 Ln5a1 Ln8a1 0.675208
Kn5an8a2 Ln5a2 Ln8a2 0.675208
Kn5an8a3 Ln5a3 Ln8a3 0.675208
Kn5an8a4 Ln5a4 Ln8a4 0.675208
Kn5an8a5 Ln5a5 Ln8a5 0.675208
Kn5an8a6 Ln5a6 Ln8a6 0.675208
Kn5an8a7 Ln5a7 Ln8a7 0.675208
Kn5an8a8 Ln5a8 Ln8a8 0.675208
Kn5anva1 Ln5a1 Lnva1 0.640637
Kn5anva2 Ln5a2 Lnva2 0.640637
Kn5anva3 Ln5a3 Lnva3 0.640637
Kn5anva4 Ln5a4 Lnva4 0.640637
Kn5anva5 Ln5a5 Lnva5 0.640637
Kn5anva6 Ln5a6 Lnva6 0.640637
Kn5anva7 Ln5a7 Lnva7 0.640637
Kn5anva8 Ln5a8 Lnva8 0.640637
Kn6an7a1 Ln6a1 Ln7a1 0.805155
Kn6an7a2 Ln6a2 Ln7a2 0.805155
Kn6an7a3 Ln6a3 Ln7a3 0.805155
Kn6an7a4 Ln6a4 Ln7a4 0.805155
Kn6an7a5 Ln6a5 Ln7a5 0.805155
Kn6an7a6 Ln6a6 Ln7a6 0.805155
Kn6an7a7 Ln6a7 Ln7a7 0.805155
Kn6an7a8 Ln6a8 Ln7a8 0.805155
Kn6an8a1 Ln6a1 Ln8a1 0.723730
Kn6an8a2 Ln6a2 Ln8a2 0.723730
Kn6an8a3 Ln6a3 Ln8a3 0.723730
Kn6an8a4 Ln6a4 Ln8a4 0.723730
Kn6an8a5 Ln6a5 Ln8a5 0.723730
Kn6an8a6 Ln6a6 Ln8a6 0.723730
Kn6an8a7 Ln6a7 Ln8a7 0.723730
Kn6an8a8 Ln6a8 Ln8a8 0.723730
Kn6anva1 Ln6a1 Lnva1 0.675208
Kn6anva2 Ln6a2 Lnva2 0.675208
Kn6anva3 Ln6a3 Lnva3 0.675208
Kn6anva4 Ln6a4 Lnva4 0.675208
Kn6anva5 Ln6a5 Lnva5 0.675208
Kn6anva6 Ln6a6 Lnva6 0.675208
Kn6anva7 Ln6a7 Lnva7 0.675208
Kn6anva8 Ln6a8 Lnva8 0.675208
Kn7an8a1 Ln7a1 Ln8a1 0.805155
Kn7an8a2 Ln7a2 Ln8a2 0.805155
Kn7an8a3 Ln7a3 Ln8a3 0.805155
Kn7an8a4 Ln7a4 Ln8a4 0.805155
Kn7an8a5 Ln7a5 Ln8a5 0.805155
Kn7an8a6 Ln7a6 Ln8a6 0.805155
Kn7an8a7 Ln7a7 Ln8a7 0.805155
Kn7an8a8 Ln7a8 Ln8a8 0.805155
Kn7anva1 Ln7a1 Lnva1 0.723730
Kn7anva2 Ln7a2 Lnva2 0.723730
Kn7anva3 Ln7a3 Lnva3 0.723730
Kn7anva4 Ln7a4 Lnva4 0.723730
Kn7anva5 Ln7a5 Lnva5 0.723730
Kn7anva6 Ln7a6 Lnva6 0.723730
Kn7anva7 Ln7a7 Lnva7 0.723730
Kn7anva8 Ln7a8 Lnva8 0.723730
Kn8anva1 Ln8a1 Lnva1 0.805155
Kn8anva2 Ln8a2 Lnva2 0.805155
Kn8anva3 Ln8a3 Lnva3 0.805155
Kn8anva4 Ln8a4 Lnva4 0.805155
Kn8anva5 Ln8a5 Lnva5 0.805155
Kn8anva6 Ln8a6 Lnva6 0.805155
Kn8anva7 Ln8a7 Lnva7 0.805155
Kn8anva8 Ln8a8 Lnva8 0.805155
Cngan1a1 TDnga1 TDn1a1 1.694350e-014
Cngan1a2 TDnga3 TDn1a3 3.388710e-014
Cngan1a3 TDnga5 TDn1a5 3.388710e-014
Cngan1a4 TDnga7 TDn1a7 3.388710e-014
Cngan1a5 TDnga9 TDn1a9 3.388710e-014
Cngan1a6 TDnga11 TDn1a11 3.388710e-014
Cngan1a7 TDnga13 TDn1a13 3.388710e-014
Cngan1a8 TDnga15 TDn1a15 3.388710e-014
Cngan1a9 TDnga17 TDn1a17 1.694350e-014
Cngan2a1 TDnga1 TDn2a1 6.546790e-015
Cngan2a2 TDnga3 TDn2a3 1.309360e-014
Cngan2a3 TDnga5 TDn2a5 1.309360e-014
Cngan2a4 TDnga7 TDn2a7 1.309360e-014
Cngan2a5 TDnga9 TDn2a9 1.309360e-014
Cngan2a6 TDnga11 TDn2a11 1.309360e-014
Cngan2a7 TDnga13 TDn2a13 1.309360e-014
Cngan2a8 TDnga15 TDn2a15 1.309360e-014
Cngan2a9 TDnga17 TDn2a17 6.546790e-015
Cngan3a1 TDnga1 TDn3a1 6.009140e-015
Cngan3a2 TDnga3 TDn3a3 1.201830e-014
Cngan3a3 TDnga5 TDn3a5 1.201830e-014
Cngan3a4 TDnga7 TDn3a7 1.201830e-014
Cngan3a5 TDnga9 TDn3a9 1.201830e-014
Cngan3a6 TDnga11 TDn3a11 1.201830e-014
Cngan3a7 TDnga13 TDn3a13 1.201830e-014
Cngan3a8 TDnga15 TDn3a15 1.201830e-014
Cngan3a9 TDnga17 TDn3a17 6.009140e-015
Cngan4a1 TDnga1 TDn4a1 5.850980e-015
Cngan4a2 TDnga3 TDn4a3 1.170200e-014
Cngan4a3 TDnga5 TDn4a5 1.170200e-014
Cngan4a4 TDnga7 TDn4a7 1.170200e-014
Cngan4a5 TDnga9 TDn4a9 1.170200e-014
Cngan4a6 TDnga11 TDn4a11 1.170200e-014
Cngan4a7 TDnga13 TDn4a13 1.170200e-014
Cngan4a8 TDnga15 TDn4a15 1.170200e-014
Cngan4a9 TDnga17 TDn4a17 5.850980e-015
Cngan5a1 TDnga1 TDn5a1 5.758530e-015
Cngan5a2 TDnga3 TDn5a3 1.151710e-014
Cngan5a3 TDnga5 TDn5a5 1.151710e-014
Cngan5a4 TDnga7 TDn5a7 1.151710e-014
Cngan5a5 TDnga9 TDn5a9 1.151710e-014
Cngan5a6 TDnga11 TDn5a11 1.151710e-014
Cngan5a7 TDnga13 TDn5a13 1.151710e-014
Cngan5a8 TDnga15 TDn5a15 1.151710e-014
Cngan5a9 TDnga17 TDn5a17 5.758530e-015
Cngan6a1 TDnga1 TDn6a1 5.724210e-015
Cngan6a2 TDnga3 TDn6a3 1.144840e-014
Cngan6a3 TDnga5 TDn6a5 1.144840e-014
Cngan6a4 TDnga7 TDn6a7 1.144840e-014
Cngan6a5 TDnga9 TDn6a9 1.144840e-014
Cngan6a6 TDnga11 TDn6a11 1.144840e-014
Cngan6a7 TDnga13 TDn6a13 1.144840e-014
Cngan6a8 TDnga15 TDn6a15 1.144840e-014
Cngan6a9 TDnga17 TDn6a17 5.724210e-015
Cngan7a1 TDnga1 TDn7a1 5.734420e-015
Cngan7a2 TDnga3 TDn7a3 1.146880e-014
Cngan7a3 TDnga5 TDn7a5 1.146880e-014
Cngan7a4 TDnga7 TDn7a7 1.146880e-014
Cngan7a5 TDnga9 TDn7a9 1.146880e-014
Cngan7a6 TDnga11 TDn7a11 1.146880e-014
Cngan7a7 TDnga13 TDn7a13 1.146880e-014
Cngan7a8 TDnga15 TDn7a15 1.146880e-014
Cngan7a9 TDnga17 TDn7a17 5.734420e-015
Cngan8a1 TDnga1 TDn8a1 5.773050e-015
Cngan8a2 TDnga3 TDn8a3 1.154610e-014
Cngan8a3 TDnga5 TDn8a5 1.154610e-014
Cngan8a4 TDnga7 TDn8a7 1.154610e-014
Cngan8a5 TDnga9 TDn8a9 1.154610e-014
Cngan8a6 TDnga11 TDn8a11 1.154610e-014
Cngan8a7 TDnga13 TDn8a13 1.154610e-014
Cngan8a8 TDnga15 TDn8a15 1.154610e-014
Cngan8a9 TDnga17 TDn8a17 5.773050e-015
Cnganva1 TDnga1 TDnva1 6.592280e-015
Cnganva2 TDnga3 TDnva3 1.318460e-014
Cnganva3 TDnga5 TDnva5 1.318460e-014
Cnganva4 TDnga7 TDnva7 1.318460e-014
Cnganva5 TDnga9 TDnva9 1.318460e-014
Cnganva6 TDnga11 TDnva11 1.318460e-014
Cnganva7 TDnga13 TDnva13 1.318460e-014
Cnganva8 TDnga15 TDnva15 1.318460e-014
Cnganva9 TDnga17 TDnva17 6.592280e-015
Cn1an2a1 TDn1a1 TDn2a1 1.586220e-014
Cn1an2a2 TDn1a3 TDn2a3 3.172450e-014
Cn1an2a3 TDn1a5 TDn2a5 3.172450e-014
Cn1an2a4 TDn1a7 TDn2a7 3.172450e-014
Cn1an2a5 TDn1a9 TDn2a9 3.172450e-014
Cn1an2a6 TDn1a11 TDn2a11 3.172450e-014
Cn1an2a7 TDn1a13 TDn2a13 3.172450e-014
Cn1an2a8 TDn1a15 TDn2a15 3.172450e-014
Cn1an2a9 TDn1a17 TDn2a17 1.586220e-014
Cn1an3a1 TDn1a1 TDn3a1 5.674250e-015
Cn1an3a2 TDn1a3 TDn3a3 1.134850e-014
Cn1an3a3 TDn1a5 TDn3a5 1.134850e-014
Cn1an3a4 TDn1a7 TDn3a7 1.134850e-014
Cn1an3a5 TDn1a9 TDn3a9 1.134850e-014
Cn1an3a6 TDn1a11 TDn3a11 1.134850e-014
Cn1an3a7 TDn1a13 TDn3a13 1.134850e-014
Cn1an3a8 TDn1a15 TDn3a15 1.134850e-014
Cn1an3a9 TDn1a17 TDn3a17 5.674250e-015
Cn1an4a1 TDn1a1 TDn4a1 5.219520e-015
Cn1an4a2 TDn1a3 TDn4a3 1.043900e-014
Cn1an4a3 TDn1a5 TDn4a5 1.043900e-014
Cn1an4a4 TDn1a7 TDn4a7 1.043900e-014
Cn1an4a5 TDn1a9 TDn4a9 1.043900e-014
Cn1an4a6 TDn1a11 TDn4a11 1.043900e-014
Cn1an4a7 TDn1a13 TDn4a13 1.043900e-014
Cn1an4a8 TDn1a15 TDn4a15 1.043900e-014
Cn1an4a9 TDn1a17 TDn4a17 5.219520e-015
Cn1an5a1 TDn1a1 TDn5a1 5.062210e-015
Cn1an5a2 TDn1a3 TDn5a3 1.012440e-014
Cn1an5a3 TDn1a5 TDn5a5 1.012440e-014
Cn1an5a4 TDn1a7 TDn5a7 1.012440e-014
Cn1an5a5 TDn1a9 TDn5a9 1.012440e-014
Cn1an5a6 TDn1a11 TDn5a11 1.012440e-014
Cn1an5a7 TDn1a13 TDn5a13 1.012440e-014
Cn1an5a8 TDn1a15 TDn5a15 1.012440e-014
Cn1an5a9 TDn1a17 TDn5a17 5.062210e-015
Cn1an6a1 TDn1a1 TDn6a1 5.003840e-015
Cn1an6a2 TDn1a3 TDn6a3 1.000770e-014
Cn1an6a3 TDn1a5 TDn6a5 1.000770e-014
Cn1an6a4 TDn1a7 TDn6a7 1.000770e-014
Cn1an6a5 TDn1a9 TDn6a9 1.000770e-014
Cn1an6a6 TDn1a11 TDn6a11 1.000770e-014
Cn1an6a7 TDn1a13 TDn6a13 1.000770e-014
Cn1an6a8 TDn1a15 TDn6a15 1.000770e-014
Cn1an6a9 TDn1a17 TDn6a17 5.003840e-015
Cn1an7a1 TDn1a1 TDn7a1 4.990870e-015
Cn1an7a2 TDn1a3 TDn7a3 9.981750e-015
Cn1an7a3 TDn1a5 TDn7a5 9.981750e-015
Cn1an7a4 TDn1a7 TDn7a7 9.981750e-015
Cn1an7a5 TDn1a9 TDn7a9 9.981750e-015
Cn1an7a6 TDn1a11 TDn7a11 9.981750e-015
Cn1an7a7 TDn1a13 TDn7a13 9.981750e-015
Cn1an7a8 TDn1a15 TDn7a15 9.981750e-015
Cn1an7a9 TDn1a17 TDn7a17 4.990870e-015
Cn1an8a1 TDn1a1 TDn8a1 5.026740e-015
Cn1an8a2 TDn1a3 TDn8a3 1.005350e-014
Cn1an8a3 TDn1a5 TDn8a5 1.005350e-014
Cn1an8a4 TDn1a7 TDn8a7 1.005350e-014
Cn1an8a5 TDn1a9 TDn8a9 1.005350e-014
Cn1an8a6 TDn1a11 TDn8a11 1.005350e-014
Cn1an8a7 TDn1a13 TDn8a13 1.005350e-014
Cn1an8a8 TDn1a15 TDn8a15 1.005350e-014
Cn1an8a9 TDn1a17 TDn8a17 5.026740e-015
Cn1anva1 TDn1a1 TDnva1 5.751040e-015
Cn1anva2 TDn1a3 TDnva3 5.751040e-015
Cn1anva3 TDn1a5 TDnva5 5.751040e-015
Cn1anva4 TDn1a7 TDnva7 5.751040e-015
Cn1anva5 TDn1a9 TDnva9 5.751040e-015
Cn1anva6 TDn1a11 TDnva11 5.751040e-015
Cn1anva7 TDn1a13 TDnva13 5.751040e-015
Cn1anva8 TDn1a15 TDnva15 5.751040e-015
Cn1anva9 TDn1a17 TDnva17 5.751040e-015
Cn2an3a1 TDn2a1 TDn3a1 1.576950e-014
Cn2an3a2 TDn2a3 TDn3a3 3.153910e-014
Cn2an3a3 TDn2a5 TDn3a5 3.153910e-014
Cn2an3a4 TDn2a7 TDn3a7 3.153910e-014
Cn2an3a5 TDn2a9 TDn3a9 3.153910e-014
Cn2an3a6 TDn2a11 TDn3a11 3.153910e-014
Cn2an3a7 TDn2a13 TDn3a13 3.153910e-014
Cn2an3a8 TDn2a15 TDn3a15 3.153910e-014
Cn2an3a9 TDn2a17 TDn3a17 1.576950e-014
Cn2an4a1 TDn2a1 TDn4a1 5.623050e-015
Cn2an4a2 TDn2a3 TDn4a3 1.124610e-014
Cn2an4a3 TDn2a5 TDn4a5 1.124610e-014
Cn2an4a4 TDn2a7 TDn4a7 1.124610e-014
Cn2an4a5 TDn2a9 TDn4a9 1.124610e-014
Cn2an4a6 TDn2a11 TDn4a11 1.124610e-014
Cn2an4a7 TDn2a13 TDn4a13 1.124610e-014
Cn2an4a8 TDn2a15 TDn4a15 1.124610e-014
Cn2an4a9 TDn2a17 TDn4a17 5.623050e-015
Cn2an5a1 TDn2a1 TDn5a1 5.149670e-015
Cn2an5a2 TDn2a3 TDn5a3 1.029930e-014
Cn2an5a3 TDn2a5 TDn5a5 1.029930e-014
Cn2an5a4 TDn2a7 TDn5a7 1.029930e-014
Cn2an5a5 TDn2a9 TDn5a9 1.029930e-014
Cn2an5a6 TDn2a11 TDn5a11 1.029930e-014
Cn2an5a7 TDn2a13 TDn5a13 1.029930e-014
Cn2an5a8 TDn2a15 TDn5a15 1.029930e-014
Cn2an5a9 TDn2a17 TDn5a17 5.149670e-015
Cn2an6a1 TDn2a1 TDn6a1 5.011480e-015
Cn2an6a2 TDn2a3 TDn6a3 1.002300e-014
Cn2an6a3 TDn2a5 TDn6a5 1.002300e-014
Cn2an6a4 TDn2a7 TDn6a7 1.002300e-014
Cn2an6a5 TDn2a9 TDn6a9 1.002300e-014
Cn2an6a6 TDn2a11 TDn6a11 1.002300e-014
Cn2an6a7 TDn2a13 TDn6a13 1.002300e-014
Cn2an6a8 TDn2a15 TDn6a15 1.002300e-014
Cn2an6a9 TDn2a17 TDn6a17 5.011480e-015
Cn2an7a1 TDn2a1 TDn7a1 4.968610e-015
Cn2an7a2 TDn2a3 TDn7a3 9.937210e-015
Cn2an7a3 TDn2a5 TDn7a5 9.937210e-015
Cn2an7a4 TDn2a7 TDn7a7 9.937210e-015
Cn2an7a5 TDn2a9 TDn7a9 9.937210e-015
Cn2an7a6 TDn2a11 TDn7a11 9.937210e-015
Cn2an7a7 TDn2a13 TDn7a13 9.937210e-015
Cn2an7a8 TDn2a15 TDn7a15 9.937210e-015
Cn2an7a9 TDn2a17 TDn7a17 4.968610e-015
Cn2an8a1 TDn2a1 TDn8a1 4.990350e-015
Cn2an8a2 TDn2a3 TDn8a3 9.980710e-015
Cn2an8a3 TDn2a5 TDn8a5 9.980710e-015
Cn2an8a4 TDn2a7 TDn8a7 9.980710e-015
Cn2an8a5 TDn2a9 TDn8a9 9.980710e-015
Cn2an8a6 TDn2a11 TDn8a11 9.980710e-015
Cn2an8a7 TDn2a13 TDn8a13 9.980710e-015
Cn2an8a8 TDn2a15 TDn8a15 9.980710e-015
Cn2an8a9 TDn2a17 TDn8a17 4.990350e-015
Cn2anva1 TDn2a1 TDnva1 5.701980e-015
Cn2anva2 TDn2a3 TDnva3 5.701980e-015
Cn2anva3 TDn2a5 TDnva5 5.701980e-015
Cn2anva4 TDn2a7 TDnva7 5.701980e-015
Cn2anva5 TDn2a9 TDnva9 5.701980e-015
Cn2anva6 TDn2a11 TDnva11 5.701980e-015
Cn2anva7 TDn2a13 TDnva13 5.701980e-015
Cn2anva8 TDn2a15 TDnva15 5.701980e-015
Cn2anva9 TDn2a17 TDnva17 5.701980e-015
Cn3an4a1 TDn3a1 TDn4a1 1.575450e-014
Cn3an4a2 TDn3a3 TDn4a3 3.150900e-014
Cn3an4a3 TDn3a5 TDn4a5 3.150900e-014
Cn3an4a4 TDn3a7 TDn4a7 3.150900e-014
Cn3an4a5 TDn3a9 TDn4a9 3.150900e-014
Cn3an4a6 TDn3a11 TDn4a11 3.150900e-014
Cn3an4a7 TDn3a13 TDn4a13 3.150900e-014
Cn3an4a8 TDn3a15 TDn4a15 3.150900e-014
Cn3an4a9 TDn3a17 TDn4a17 1.575450e-014
Cn3an5a1 TDn3a1 TDn5a1 5.588630e-015
Cn3an5a2 TDn3a3 TDn5a3 1.117730e-014
Cn3an5a3 TDn3a5 TDn5a5 1.117730e-014
Cn3an5a4 TDn3a7 TDn5a7 1.117730e-014
Cn3an5a5 TDn3a9 TDn5a9 1.117730e-014
Cn3an5a6 TDn3a11 TDn5a11 1.117730e-014
Cn3an5a7 TDn3a13 TDn5a13 1.117730e-014
Cn3an5a8 TDn3a15 TDn5a15 1.117730e-014
Cn3an5a9 TDn3a17 TDn5a17 5.588630e-015
Cn3an6a1 TDn3a1 TDn6a1 5.135110e-015
Cn3an6a2 TDn3a3 TDn6a3 1.027020e-014
Cn3an6a3 TDn3a5 TDn6a5 1.027020e-014
Cn3an6a4 TDn3a7 TDn6a7 1.027020e-014
Cn3an6a5 TDn3a9 TDn6a9 1.027020e-014
Cn3an6a6 TDn3a11 TDn6a11 1.027020e-014
Cn3an6a7 TDn3a13 TDn6a13 1.027020e-014
Cn3an6a8 TDn3a15 TDn6a15 1.027020e-014
Cn3an6a9 TDn3a17 TDn6a17 5.135110e-015
Cn3an7a1 TDn3a1 TDn7a1 5.012180e-015
Cn3an7a2 TDn3a3 TDn7a3 1.002440e-014
Cn3an7a3 TDn3a5 TDn7a5 1.002440e-014
Cn3an7a4 TDn3a7 TDn7a7 1.002440e-014
Cn3an7a5 TDn3a9 TDn7a9 1.002440e-014
Cn3an7a6 TDn3a11 TDn7a11 1.002440e-014
Cn3an7a7 TDn3a13 TDn7a13 1.002440e-014
Cn3an7a8 TDn3a15 TDn7a15 1.002440e-014
Cn3an7a9 TDn3a17 TDn7a17 5.012180e-015
Cn3an8a1 TDn3a1 TDn8a1 5.004030e-015
Cn3an8a2 TDn3a3 TDn8a3 1.000810e-014
Cn3an8a3 TDn3a5 TDn8a5 1.000810e-014
Cn3an8a4 TDn3a7 TDn8a7 1.000810e-014
Cn3an8a5 TDn3a9 TDn8a9 1.000810e-014
Cn3an8a6 TDn3a11 TDn8a11 1.000810e-014
Cn3an8a7 TDn3a13 TDn8a13 1.000810e-014
Cn3an8a8 TDn3a15 TDn8a15 1.000810e-014
Cn3an8a9 TDn3a17 TDn8a17 5.004030e-015
Cn3anva1 TDn3a1 TDnva1 5.703560e-015
Cn3anva2 TDn3a3 TDnva3 5.703560e-015
Cn3anva3 TDn3a5 TDnva5 5.703560e-015
Cn3anva4 TDn3a7 TDnva7 5.703560e-015
Cn3anva5 TDn3a9 TDnva9 5.703560e-015
Cn3anva6 TDn3a11 TDnva11 5.703560e-015
Cn3anva7 TDn3a13 TDnva13 5.703560e-015
Cn3anva8 TDn3a15 TDnva15 5.703560e-015
Cn3anva9 TDn3a17 TDnva17 5.703560e-015
Cn4an5a1 TDn4a1 TDn5a1 1.573240e-014
Cn4an5a2 TDn4a3 TDn5a3 3.146480e-014
Cn4an5a3 TDn4a5 TDn5a5 3.146480e-014
Cn4an5a4 TDn4a7 TDn5a7 3.146480e-014
Cn4an5a5 TDn4a9 TDn5a9 3.146480e-014
Cn4an5a6 TDn4a11 TDn5a11 3.146480e-014
Cn4an5a7 TDn4a13 TDn5a13 3.146480e-014
Cn4an5a8 TDn4a15 TDn5a15 3.146480e-014
Cn4an5a9 TDn4a17 TDn5a17 1.573240e-014
Cn4an6a1 TDn4a1 TDn6a1 5.586810e-015
Cn4an6a2 TDn4a3 TDn6a3 1.117360e-014
Cn4an6a3 TDn4a5 TDn6a5 1.117360e-014
Cn4an6a4 TDn4a7 TDn6a7 1.117360e-014
Cn4an6a5 TDn4a9 TDn6a9 1.117360e-014
Cn4an6a6 TDn4a11 TDn6a11 1.117360e-014
Cn4an6a7 TDn4a13 TDn6a13 1.117360e-014
Cn4an6a8 TDn4a15 TDn6a15 1.117360e-014
Cn4an6a9 TDn4a17 TDn6a17 5.586810e-015
Cn4an7a1 TDn4a1 TDn7a1 5.148610e-015
Cn4an7a2 TDn4a3 TDn7a3 1.029720e-014
Cn4an7a3 TDn4a5 TDn7a5 1.029720e-014
Cn4an7a4 TDn4a7 TDn7a7 1.029720e-014
Cn4an7a5 TDn4a9 TDn7a9 1.029720e-014
Cn4an7a6 TDn4a11 TDn7a11 1.029720e-014
Cn4an7a7 TDn4a13 TDn7a13 1.029720e-014
Cn4an7a8 TDn4a15 TDn7a15 1.029720e-014
Cn4an7a9 TDn4a17 TDn7a17 5.148610e-015
Cn4an8a1 TDn4a1 TDn8a1 5.060570e-015
Cn4an8a2 TDn4a3 TDn8a3 1.012110e-014
Cn4an8a3 TDn4a5 TDn8a5 1.012110e-014
Cn4an8a4 TDn4a7 TDn8a7 1.012110e-014
Cn4an8a5 TDn4a9 TDn8a9 1.012110e-014
Cn4an8a6 TDn4a11 TDn8a11 1.012110e-014
Cn4an8a7 TDn4a13 TDn8a13 1.012110e-014
Cn4an8a8 TDn4a15 TDn8a15 1.012110e-014
Cn4an8a9 TDn4a17 TDn8a17 5.060570e-015
Cn4anva1 TDn4a1 TDnva1 5.736010e-015
Cn4anva2 TDn4a3 TDnva3 5.736010e-015
Cn4anva3 TDn4a5 TDnva5 5.736010e-015
Cn4anva4 TDn4a7 TDnva7 5.736010e-015
Cn4anva5 TDn4a9 TDnva9 5.736010e-015
Cn4anva6 TDn4a11 TDnva11 5.736010e-015
Cn4anva7 TDn4a13 TDnva13 5.736010e-015
Cn4anva8 TDn4a15 TDnva15 5.736010e-015
Cn4anva9 TDn4a17 TDnva17 5.736010e-015
Cn5an6a1 TDn5a1 TDn6a1 1.575710e-014
Cn5an6a2 TDn5a3 TDn6a3 3.151420e-014
Cn5an6a3 TDn5a5 TDn6a5 3.151420e-014
Cn5an6a4 TDn5a7 TDn6a7 3.151420e-014
Cn5an6a5 TDn5a9 TDn6a9 3.151420e-014
Cn5an6a6 TDn5a11 TDn6a11 3.151420e-014
Cn5an6a7 TDn5a13 TDn6a13 3.151420e-014
Cn5an6a8 TDn5a15 TDn6a15 3.151420e-014
Cn5an6a9 TDn5a17 TDn6a17 1.575710e-014
Cn5an7a1 TDn5a1 TDn7a1 5.608560e-015
Cn5an7a2 TDn5a3 TDn7a3 1.121710e-014
Cn5an7a3 TDn5a5 TDn7a5 1.121710e-014
Cn5an7a4 TDn5a7 TDn7a7 1.121710e-014
Cn5an7a5 TDn5a9 TDn7a9 1.121710e-014
Cn5an7a6 TDn5a11 TDn7a11 1.121710e-014
Cn5an7a7 TDn5a13 TDn7a13 1.121710e-014
Cn5an7a8 TDn5a15 TDn7a15 1.121710e-014
Cn5an7a9 TDn5a17 TDn7a17 5.608560e-015
Cn5an8a1 TDn5a1 TDn8a1 5.204690e-015
Cn5an8a2 TDn5a3 TDn8a3 1.040940e-014
Cn5an8a3 TDn5a5 TDn8a5 1.040940e-014
Cn5an8a4 TDn5a7 TDn8a7 1.040940e-014
Cn5an8a5 TDn5a9 TDn8a9 1.040940e-014
Cn5an8a6 TDn5a11 TDn8a11 1.040940e-014
Cn5an8a7 TDn5a13 TDn8a13 1.040940e-014
Cn5an8a8 TDn5a15 TDn8a15 1.040940e-014
Cn5an8a9 TDn5a17 TDn8a17 5.204690e-015
Cn5anva1 TDn5a1 TDnva1 5.818520e-015
Cn5anva2 TDn5a3 TDnva3 5.818520e-015
Cn5anva3 TDn5a5 TDnva5 5.818520e-015
Cn5anva4 TDn5a7 TDnva7 5.818520e-015
Cn5anva5 TDn5a9 TDnva9 5.818520e-015
Cn5anva6 TDn5a11 TDnva11 5.818520e-015
Cn5anva7 TDn5a13 TDnva13 5.818520e-015
Cn5anva8 TDn5a15 TDnva15 5.818520e-015
Cn5anva9 TDn5a17 TDnva17 5.818520e-015
Cn6an7a1 TDn6a1 TDn7a1 1.578870e-014
Cn6an7a2 TDn6a3 TDn7a3 3.157750e-014
Cn6an7a3 TDn6a5 TDn7a5 3.157750e-014
Cn6an7a4 TDn6a7 TDn7a7 3.157750e-014
Cn6an7a5 TDn6a9 TDn7a9 3.157750e-014
Cn6an7a6 TDn6a11 TDn7a11 3.157750e-014
Cn6an7a7 TDn6a13 TDn7a13 3.157750e-014
Cn6an7a8 TDn6a15 TDn7a15 3.157750e-014
Cn6an7a9 TDn6a17 TDn7a17 1.578870e-014
Cn6an8a1 TDn6a1 TDn8a1 5.673080e-015
Cn6an8a2 TDn6a3 TDn8a3 1.134620e-014
Cn6an8a3 TDn6a5 TDn8a5 1.134620e-014
Cn6an8a4 TDn6a7 TDn8a7 1.134620e-014
Cn6an8a5 TDn6a9 TDn8a9 1.134620e-014
Cn6an8a6 TDn6a11 TDn8a11 1.134620e-014
Cn6an8a7 TDn6a13 TDn8a13 1.134620e-014
Cn6an8a8 TDn6a15 TDn8a15 1.134620e-014
Cn6an8a9 TDn6a17 TDn8a17 5.673080e-015
Cn6anva1 TDn6a1 TDnva1 6.001130e-015
Cn6anva2 TDn6a3 TDnva3 6.001130e-015
Cn6anva3 TDn6a5 TDnva5 6.001130e-015
Cn6anva4 TDn6a7 TDnva7 6.001130e-015
Cn6anva5 TDn6a9 TDnva9 6.001130e-015
Cn6anva6 TDn6a11 TDnva11 6.001130e-015
Cn6anva7 TDn6a13 TDnva13 6.001130e-015
Cn6anva8 TDn6a15 TDnva15 6.001130e-015
Cn6anva9 TDn6a17 TDnva17 6.001130e-015
Cn7an8a1 TDn7a1 TDn8a1 1.587490e-014
Cn7an8a2 TDn7a3 TDn8a3 3.174970e-014
Cn7an8a3 TDn7a5 TDn8a5 3.174970e-014
Cn7an8a4 TDn7a7 TDn8a7 3.174970e-014
Cn7an8a5 TDn7a9 TDn8a9 3.174970e-014
Cn7an8a6 TDn7a11 TDn8a11 3.174970e-014
Cn7an8a7 TDn7a13 TDn8a13 3.174970e-014
Cn7an8a8 TDn7a15 TDn8a15 3.174970e-014
Cn7an8a9 TDn7a17 TDn8a17 1.587490e-014
Cn7anva1 TDn7a1 TDnva1 6.511580e-015
Cn7anva2 TDn7a3 TDnva3 6.511580e-015
Cn7anva3 TDn7a5 TDnva5 6.511580e-015
Cn7anva4 TDn7a7 TDnva7 6.511580e-015
Cn7anva5 TDn7a9 TDnva9 6.511580e-015
Cn7anva6 TDn7a11 TDnva11 6.511580e-015
Cn7anva7 TDn7a13 TDnva13 6.511580e-015
Cn7anva8 TDn7a15 TDnva15 6.511580e-015
Cn7anva9 TDn7a17 TDnva17 6.511580e-015
Cn8anva1 TDn8a1 TDnva1 1.690880e-014
Cn8anva2 TDn8a3 TDnva3 1.690880e-014
Cn8anva3 TDn8a5 TDnva5 1.690880e-014
Cn8anva4 TDn8a7 TDnva7 1.690880e-014
Cn8anva5 TDn8a9 TDnva9 1.690880e-014
Cn8anva6 TDn8a11 TDnva11 1.690880e-014
Cn8anva7 TDn8a13 TDnva13 1.690880e-014
Cn8anva8 TDn8a15 TDnva15 1.690880e-014
Cn8anva9 TDn8a17 TDnva17 1.690880e-014
.ENDS intercon
*.output v<cout1>
*.op 
*.AC LIN 1000 0 10G 
.Tran 1e-12 1e-9 
.probe  V(TDn1a9)  V(TDn2a9)  V(TDn3a9)  V(TDn4a9)  V(TDn5a9)  V(TDn6a9)  V(TDn7a9)  V(TDn8a9)  V(TDn8a1)  V(TDn7a1)  V(TDn6a1)  V(TDn5a1)  V(TDn4a1)  V(TDn3a1)  V(TDn2a1)  V(TDn1a1) 
.print  V(TDn1a9)  V(TDn2a9)  V(TDn3a9)  V(TDn4a9)  V(TDn5a9)  V(TDn6a9)  V(TDn7a9)  V(TDn8a9)  V(TDn8a1)  V(TDn7a1)  V(TDn6a1)  V(TDn5a1)  V(TDn4a1)  V(TDn3a1)  V(TDn2a1)  V(TDn1a1) 
.end
