*A distribution linear circuit for line 14 segment 16.
Vin1 TDvn1a1 0 AC 1

Rin1 TDvn1a1 TDn1a1 10

Rs2 TDvn2a1 0 0.1
Rs3 TDvn3a1 0 0.1
Rs4 TDvn4a1 0 0.1
Rs5 TDvn5a1 0 0.1
Rs6 TDvn6a1 0 0.1
Rs7 TDvn7a1 0 0.1
Rs8 TDvn8a1 0 0.1
Rs9 TDvn9a1 0 0.1
Rs10 TDvn10a1 0 0.1
Rs11 TDvn11a1 0 0.1
Rs12 TDvn12a1 0 0.1

Rgndg TDnga1 0 1
Rgnd2 TDn2a1 0 10
Rgnd3 TDn3a1 0 10
Rgnd4 TDn4a1 0 10
Rgnd5 TDn5a1 0 10
Rgnd6 TDn6a1 0 10
Rgnd7 TDn7a1 0 10
Rgnd8 TDn8a1 0 10
Rgnd9 TDn9a1 0 10
Rgnd10 TDn10a1 0 10
Rgnd11 TDn11a1 0 10
Rgnd12 TDn12a1 0 10
Rgndv TDnva1 0 1

RRR TDnga9 TDnva9 1
Cout1 TDn1a9 TDnga9 0.1p
Cout2 TDn2a9 TDnga9 0.1p
Cout3 TDn3a9 TDnga9 0.1p
Cout4 TDn4a9 TDnga9 0.1p
Cout5 TDn5a9 TDnga9 0.1p
Cout6 TDn6a9 TDnga9 0.1p
Cout7 TDn7a9 TDnga9 0.1p
Cout8 TDn8a9 TDnga9 0.1p
Cout9 TDn9a9 TDnga9 0.1p
Cout10 TDn10a9 TDnga9 0.1p
Cout11 TDn11a9 TDnga9 0.1p
Cout12 TDn12a9 TDnga9 0.1p

X1 TDnga1 TDnga9 TDn1a1 TDn1a9 TDn2a1 TDn2a9 TDn3a1 TDn3a9 TDn4a1 TDn4a9 TDn5a1 TDn5a9 TDn6a1 TDn6a9 TDn7a1 TDn7a9 TDn8a1 TDn8a9 TDn9a1 TDn9a9 TDn10a1 TDn10a9 TDn11a1 TDn11a9 TDn12a1 TDn12a9 TDnva1 TDnva9 intercon
.SUBCKT intercon TDnga1 TDnga33 TDn1a1 TDn1a33 TDn2a1 TDn2a33 TDn3a1 TDn3a33 TDn4a1 TDn4a33 TDn5a1 TDn5a33 TDn6a1 TDn6a33 TDn7a1 TDn7a33 TDn8a1 TDn8a33 TDn9a1 TDn9a33 TDn10a1 TDn10a33 TDn11a1 TDn11a33 TDn12a1 TDn12a33 TDnva1 TDnva33

Rnga1 TDnga1 TDnga2 2
Rnga2 TDnga3 TDnga4 2
Rnga3 TDnga5 TDnga6 2
Rnga4 TDnga7 TDnga8 2
Rnga5 TDnga9 TDnga10 2
Rnga6 TDnga11 TDnga12 2
Rnga7 TDnga13 TDnga14 2
Rnga8 TDnga15 TDnga16 2
Rnga9 TDnga17 TDnga18 2
Rnga10 TDnga19 TDnga20 2
Rnga11 TDnga21 TDnga22 2
Rnga12 TDnga23 TDnga24 2
Rnga13 TDnga25 TDnga26 2
Rnga14 TDnga27 TDnga28 2
Rnga15 TDnga29 TDnga30 2
Rnga16 TDnga31 TDnga32 2
Rn1a1 TDn1a1 TDn1a2 2
Rn1a2 TDn1a3 TDn1a4 2
Rn1a3 TDn1a5 TDn1a6 2
Rn1a4 TDn1a7 TDn1a8 2
Rn1a5 TDn1a9 TDn1a10 2
Rn1a6 TDn1a11 TDn1a12 2
Rn1a7 TDn1a13 TDn1a14 2
Rn1a8 TDn1a15 TDn1a16 2
Rn1a9 TDn1a17 TDn1a18 2
Rn1a10 TDn1a19 TDn1a20 2
Rn1a11 TDn1a21 TDn1a22 2
Rn1a12 TDn1a23 TDn1a24 2
Rn1a13 TDn1a25 TDn1a26 2
Rn1a14 TDn1a27 TDn1a28 2
Rn1a15 TDn1a29 TDn1a30 2
Rn1a16 TDn1a31 TDn1a32 2
Rn2a1 TDn2a1 TDn2a2 2
Rn2a2 TDn2a3 TDn2a4 2
Rn2a3 TDn2a5 TDn2a6 2
Rn2a4 TDn2a7 TDn2a8 2
Rn2a5 TDn2a9 TDn2a10 2
Rn2a6 TDn2a11 TDn2a12 2
Rn2a7 TDn2a13 TDn2a14 2
Rn2a8 TDn2a15 TDn2a16 2
Rn2a9 TDn2a17 TDn2a18 2
Rn2a10 TDn2a19 TDn2a20 2
Rn2a11 TDn2a21 TDn2a22 2
Rn2a12 TDn2a23 TDn2a24 2
Rn2a13 TDn2a25 TDn2a26 2
Rn2a14 TDn2a27 TDn2a28 2
Rn2a15 TDn2a29 TDn2a30 2
Rn2a16 TDn2a31 TDn2a32 2
Rn3a1 TDn3a1 TDn3a2 2
Rn3a2 TDn3a3 TDn3a4 2
Rn3a3 TDn3a5 TDn3a6 2
Rn3a4 TDn3a7 TDn3a8 2
Rn3a5 TDn3a9 TDn3a10 2
Rn3a6 TDn3a11 TDn3a12 2
Rn3a7 TDn3a13 TDn3a14 2
Rn3a8 TDn3a15 TDn3a16 2
Rn3a9 TDn3a17 TDn3a18 2
Rn3a10 TDn3a19 TDn3a20 2
Rn3a11 TDn3a21 TDn3a22 2
Rn3a12 TDn3a23 TDn3a24 2
Rn3a13 TDn3a25 TDn3a26 2
Rn3a14 TDn3a27 TDn3a28 2
Rn3a15 TDn3a29 TDn3a30 2
Rn3a16 TDn3a31 TDn3a32 2
Rn4a1 TDn4a1 TDn4a2 2
Rn4a2 TDn4a3 TDn4a4 2
Rn4a3 TDn4a5 TDn4a6 2
Rn4a4 TDn4a7 TDn4a8 2
Rn4a5 TDn4a9 TDn4a10 2
Rn4a6 TDn4a11 TDn4a12 2
Rn4a7 TDn4a13 TDn4a14 2
Rn4a8 TDn4a15 TDn4a16 2
Rn4a9 TDn4a17 TDn4a18 2
Rn4a10 TDn4a19 TDn4a20 2
Rn4a11 TDn4a21 TDn4a22 2
Rn4a12 TDn4a23 TDn4a24 2
Rn4a13 TDn4a25 TDn4a26 2
Rn4a14 TDn4a27 TDn4a28 2
Rn4a15 TDn4a29 TDn4a30 2
Rn4a16 TDn4a31 TDn4a32 2
Rn5a1 TDn5a1 TDn5a2 2
Rn5a2 TDn5a3 TDn5a4 2
Rn5a3 TDn5a5 TDn5a6 2
Rn5a4 TDn5a7 TDn5a8 2
Rn5a5 TDn5a9 TDn5a10 2
Rn5a6 TDn5a11 TDn5a12 2
Rn5a7 TDn5a13 TDn5a14 2
Rn5a8 TDn5a15 TDn5a16 2
Rn5a9 TDn5a17 TDn5a18 2
Rn5a10 TDn5a19 TDn5a20 2
Rn5a11 TDn5a21 TDn5a22 2
Rn5a12 TDn5a23 TDn5a24 2
Rn5a13 TDn5a25 TDn5a26 2
Rn5a14 TDn5a27 TDn5a28 2
Rn5a15 TDn5a29 TDn5a30 2
Rn5a16 TDn5a31 TDn5a32 2
Rn6a1 TDn6a1 TDn6a2 2
Rn6a2 TDn6a3 TDn6a4 2
Rn6a3 TDn6a5 TDn6a6 2
Rn6a4 TDn6a7 TDn6a8 2
Rn6a5 TDn6a9 TDn6a10 2
Rn6a6 TDn6a11 TDn6a12 2
Rn6a7 TDn6a13 TDn6a14 2
Rn6a8 TDn6a15 TDn6a16 2
Rn6a9 TDn6a17 TDn6a18 2
Rn6a10 TDn6a19 TDn6a20 2
Rn6a11 TDn6a21 TDn6a22 2
Rn6a12 TDn6a23 TDn6a24 2
Rn6a13 TDn6a25 TDn6a26 2
Rn6a14 TDn6a27 TDn6a28 2
Rn6a15 TDn6a29 TDn6a30 2
Rn6a16 TDn6a31 TDn6a32 2
Rn7a1 TDn7a1 TDn7a2 2
Rn7a2 TDn7a3 TDn7a4 2
Rn7a3 TDn7a5 TDn7a6 2
Rn7a4 TDn7a7 TDn7a8 2
Rn7a5 TDn7a9 TDn7a10 2
Rn7a6 TDn7a11 TDn7a12 2
Rn7a7 TDn7a13 TDn7a14 2
Rn7a8 TDn7a15 TDn7a16 2
Rn7a9 TDn7a17 TDn7a18 2
Rn7a10 TDn7a19 TDn7a20 2
Rn7a11 TDn7a21 TDn7a22 2
Rn7a12 TDn7a23 TDn7a24 2
Rn7a13 TDn7a25 TDn7a26 2
Rn7a14 TDn7a27 TDn7a28 2
Rn7a15 TDn7a29 TDn7a30 2
Rn7a16 TDn7a31 TDn7a32 2
Rn8a1 TDn8a1 TDn8a2 2
Rn8a2 TDn8a3 TDn8a4 2
Rn8a3 TDn8a5 TDn8a6 2
Rn8a4 TDn8a7 TDn8a8 2
Rn8a5 TDn8a9 TDn8a10 2
Rn8a6 TDn8a11 TDn8a12 2
Rn8a7 TDn8a13 TDn8a14 2
Rn8a8 TDn8a15 TDn8a16 2
Rn8a9 TDn8a17 TDn8a18 2
Rn8a10 TDn8a19 TDn8a20 2
Rn8a11 TDn8a21 TDn8a22 2
Rn8a12 TDn8a23 TDn8a24 2
Rn8a13 TDn8a25 TDn8a26 2
Rn8a14 TDn8a27 TDn8a28 2
Rn8a15 TDn8a29 TDn8a30 2
Rn8a16 TDn8a31 TDn8a32 2
Rn9a1 TDn9a1 TDn9a2 2
Rn9a2 TDn9a3 TDn9a4 2
Rn9a3 TDn9a5 TDn9a6 2
Rn9a4 TDn9a7 TDn9a8 2
Rn9a5 TDn9a9 TDn9a10 2
Rn9a6 TDn9a11 TDn9a12 2
Rn9a7 TDn9a13 TDn9a14 2
Rn9a8 TDn9a15 TDn9a16 2
Rn9a9 TDn9a17 TDn9a18 2
Rn9a10 TDn9a19 TDn9a20 2
Rn9a11 TDn9a21 TDn9a22 2
Rn9a12 TDn9a23 TDn9a24 2
Rn9a13 TDn9a25 TDn9a26 2
Rn9a14 TDn9a27 TDn9a28 2
Rn9a15 TDn9a29 TDn9a30 2
Rn9a16 TDn9a31 TDn9a32 2
Rn10a1 TDn10a1 TDn10a2 2
Rn10a2 TDn10a3 TDn10a4 2
Rn10a3 TDn10a5 TDn10a6 2
Rn10a4 TDn10a7 TDn10a8 2
Rn10a5 TDn10a9 TDn10a10 2
Rn10a6 TDn10a11 TDn10a12 2
Rn10a7 TDn10a13 TDn10a14 2
Rn10a8 TDn10a15 TDn10a16 2
Rn10a9 TDn10a17 TDn10a18 2
Rn10a10 TDn10a19 TDn10a20 2
Rn10a11 TDn10a21 TDn10a22 2
Rn10a12 TDn10a23 TDn10a24 2
Rn10a13 TDn10a25 TDn10a26 2
Rn10a14 TDn10a27 TDn10a28 2
Rn10a15 TDn10a29 TDn10a30 2
Rn10a16 TDn10a31 TDn10a32 2
Rn11a1 TDn11a1 TDn11a2 2
Rn11a2 TDn11a3 TDn11a4 2
Rn11a3 TDn11a5 TDn11a6 2
Rn11a4 TDn11a7 TDn11a8 2
Rn11a5 TDn11a9 TDn11a10 2
Rn11a6 TDn11a11 TDn11a12 2
Rn11a7 TDn11a13 TDn11a14 2
Rn11a8 TDn11a15 TDn11a16 2
Rn11a9 TDn11a17 TDn11a18 2
Rn11a10 TDn11a19 TDn11a20 2
Rn11a11 TDn11a21 TDn11a22 2
Rn11a12 TDn11a23 TDn11a24 2
Rn11a13 TDn11a25 TDn11a26 2
Rn11a14 TDn11a27 TDn11a28 2
Rn11a15 TDn11a29 TDn11a30 2
Rn11a16 TDn11a31 TDn11a32 2
Rn12a1 TDn12a1 TDn12a2 2
Rn12a2 TDn12a3 TDn12a4 2
Rn12a3 TDn12a5 TDn12a6 2
Rn12a4 TDn12a7 TDn12a8 2
Rn12a5 TDn12a9 TDn12a10 2
Rn12a6 TDn12a11 TDn12a12 2
Rn12a7 TDn12a13 TDn12a14 2
Rn12a8 TDn12a15 TDn12a16 2
Rn12a9 TDn12a17 TDn12a18 2
Rn12a10 TDn12a19 TDn12a20 2
Rn12a11 TDn12a21 TDn12a22 2
Rn12a12 TDn12a23 TDn12a24 2
Rn12a13 TDn12a25 TDn12a26 2
Rn12a14 TDn12a27 TDn12a28 2
Rn12a15 TDn12a29 TDn12a30 2
Rn12a16 TDn12a31 TDn12a32 2
Rnva1 TDnva1 TDnva2 2
Rnva2 TDnva3 TDnva4 2
Rnva3 TDnva5 TDnva6 2
Rnva4 TDnva7 TDnva8 2
Rnva5 TDnva9 TDnva10 2
Rnva6 TDnva11 TDnva12 2
Rnva7 TDnva13 TDnva14 2
Rnva8 TDnva15 TDnva16 2
Rnva9 TDnva17 TDnva18 2
Rnva10 TDnva19 TDnva20 2
Rnva11 TDnva21 TDnva22 2
Rnva12 TDnva23 TDnva24 2
Rnva13 TDnva25 TDnva26 2
Rnva14 TDnva27 TDnva28 2
Rnva15 TDnva29 TDnva30 2
Rnva16 TDnva31 TDnva32 2
Lnga1 TDnga2 TDnga3 1e-9
Lnga2 TDnga4 TDnga5 1e-9
Lnga3 TDnga6 TDnga7 1e-9
Lnga4 TDnga8 TDnga9 1e-9
Lnga5 TDnga10 TDnga11 1e-9
Lnga6 TDnga12 TDnga13 1e-9
Lnga7 TDnga14 TDnga15 1e-9
Lnga8 TDnga16 TDnga17 1e-9
Lnga9 TDnga18 TDnga19 1e-9
Lnga10 TDnga20 TDnga21 1e-9
Lnga11 TDnga22 TDnga23 1e-9
Lnga12 TDnga24 TDnga25 1e-9
Lnga13 TDnga26 TDnga27 1e-9
Lnga14 TDnga28 TDnga29 1e-9
Lnga15 TDnga30 TDnga31 1e-9
Lnga16 TDnga32 TDnga33 1e-9
Ln1a1 TDn1a2 TDn1a3 1e-9
Ln1a2 TDn1a4 TDn1a5 1e-9
Ln1a3 TDn1a6 TDn1a7 1e-9
Ln1a4 TDn1a8 TDn1a9 1e-9
Ln1a5 TDn1a10 TDn1a11 1e-9
Ln1a6 TDn1a12 TDn1a13 1e-9
Ln1a7 TDn1a14 TDn1a15 1e-9
Ln1a8 TDn1a16 TDn1a17 1e-9
Ln1a9 TDn1a18 TDn1a19 1e-9
Ln1a10 TDn1a20 TDn1a21 1e-9
Ln1a11 TDn1a22 TDn1a23 1e-9
Ln1a12 TDn1a24 TDn1a25 1e-9
Ln1a13 TDn1a26 TDn1a27 1e-9
Ln1a14 TDn1a28 TDn1a29 1e-9
Ln1a15 TDn1a30 TDn1a31 1e-9
Ln1a16 TDn1a32 TDn1a33 1e-9
Ln2a1 TDn2a2 TDn2a3 1e-9
Ln2a2 TDn2a4 TDn2a5 1e-9
Ln2a3 TDn2a6 TDn2a7 1e-9
Ln2a4 TDn2a8 TDn2a9 1e-9
Ln2a5 TDn2a10 TDn2a11 1e-9
Ln2a6 TDn2a12 TDn2a13 1e-9
Ln2a7 TDn2a14 TDn2a15 1e-9
Ln2a8 TDn2a16 TDn2a17 1e-9
Ln2a9 TDn2a18 TDn2a19 1e-9
Ln2a10 TDn2a20 TDn2a21 1e-9
Ln2a11 TDn2a22 TDn2a23 1e-9
Ln2a12 TDn2a24 TDn2a25 1e-9
Ln2a13 TDn2a26 TDn2a27 1e-9
Ln2a14 TDn2a28 TDn2a29 1e-9
Ln2a15 TDn2a30 TDn2a31 1e-9
Ln2a16 TDn2a32 TDn2a33 1e-9
Ln3a1 TDn3a2 TDn3a3 1e-9
Ln3a2 TDn3a4 TDn3a5 1e-9
Ln3a3 TDn3a6 TDn3a7 1e-9
Ln3a4 TDn3a8 TDn3a9 1e-9
Ln3a5 TDn3a10 TDn3a11 1e-9
Ln3a6 TDn3a12 TDn3a13 1e-9
Ln3a7 TDn3a14 TDn3a15 1e-9
Ln3a8 TDn3a16 TDn3a17 1e-9
Ln3a9 TDn3a18 TDn3a19 1e-9
Ln3a10 TDn3a20 TDn3a21 1e-9
Ln3a11 TDn3a22 TDn3a23 1e-9
Ln3a12 TDn3a24 TDn3a25 1e-9
Ln3a13 TDn3a26 TDn3a27 1e-9
Ln3a14 TDn3a28 TDn3a29 1e-9
Ln3a15 TDn3a30 TDn3a31 1e-9
Ln3a16 TDn3a32 TDn3a33 1e-9
Ln4a1 TDn4a2 TDn4a3 1e-9
Ln4a2 TDn4a4 TDn4a5 1e-9
Ln4a3 TDn4a6 TDn4a7 1e-9
Ln4a4 TDn4a8 TDn4a9 1e-9
Ln4a5 TDn4a10 TDn4a11 1e-9
Ln4a6 TDn4a12 TDn4a13 1e-9
Ln4a7 TDn4a14 TDn4a15 1e-9
Ln4a8 TDn4a16 TDn4a17 1e-9
Ln4a9 TDn4a18 TDn4a19 1e-9
Ln4a10 TDn4a20 TDn4a21 1e-9
Ln4a11 TDn4a22 TDn4a23 1e-9
Ln4a12 TDn4a24 TDn4a25 1e-9
Ln4a13 TDn4a26 TDn4a27 1e-9
Ln4a14 TDn4a28 TDn4a29 1e-9
Ln4a15 TDn4a30 TDn4a31 1e-9
Ln4a16 TDn4a32 TDn4a33 1e-9
Ln5a1 TDn5a2 TDn5a3 1e-9
Ln5a2 TDn5a4 TDn5a5 1e-9
Ln5a3 TDn5a6 TDn5a7 1e-9
Ln5a4 TDn5a8 TDn5a9 1e-9
Ln5a5 TDn5a10 TDn5a11 1e-9
Ln5a6 TDn5a12 TDn5a13 1e-9
Ln5a7 TDn5a14 TDn5a15 1e-9
Ln5a8 TDn5a16 TDn5a17 1e-9
Ln5a9 TDn5a18 TDn5a19 1e-9
Ln5a10 TDn5a20 TDn5a21 1e-9
Ln5a11 TDn5a22 TDn5a23 1e-9
Ln5a12 TDn5a24 TDn5a25 1e-9
Ln5a13 TDn5a26 TDn5a27 1e-9
Ln5a14 TDn5a28 TDn5a29 1e-9
Ln5a15 TDn5a30 TDn5a31 1e-9
Ln5a16 TDn5a32 TDn5a33 1e-9
Ln6a1 TDn6a2 TDn6a3 1e-9
Ln6a2 TDn6a4 TDn6a5 1e-9
Ln6a3 TDn6a6 TDn6a7 1e-9
Ln6a4 TDn6a8 TDn6a9 1e-9
Ln6a5 TDn6a10 TDn6a11 1e-9
Ln6a6 TDn6a12 TDn6a13 1e-9
Ln6a7 TDn6a14 TDn6a15 1e-9
Ln6a8 TDn6a16 TDn6a17 1e-9
Ln6a9 TDn6a18 TDn6a19 1e-9
Ln6a10 TDn6a20 TDn6a21 1e-9
Ln6a11 TDn6a22 TDn6a23 1e-9
Ln6a12 TDn6a24 TDn6a25 1e-9
Ln6a13 TDn6a26 TDn6a27 1e-9
Ln6a14 TDn6a28 TDn6a29 1e-9
Ln6a15 TDn6a30 TDn6a31 1e-9
Ln6a16 TDn6a32 TDn6a33 1e-9
Ln7a1 TDn7a2 TDn7a3 1e-9
Ln7a2 TDn7a4 TDn7a5 1e-9
Ln7a3 TDn7a6 TDn7a7 1e-9
Ln7a4 TDn7a8 TDn7a9 1e-9
Ln7a5 TDn7a10 TDn7a11 1e-9
Ln7a6 TDn7a12 TDn7a13 1e-9
Ln7a7 TDn7a14 TDn7a15 1e-9
Ln7a8 TDn7a16 TDn7a17 1e-9
Ln7a9 TDn7a18 TDn7a19 1e-9
Ln7a10 TDn7a20 TDn7a21 1e-9
Ln7a11 TDn7a22 TDn7a23 1e-9
Ln7a12 TDn7a24 TDn7a25 1e-9
Ln7a13 TDn7a26 TDn7a27 1e-9
Ln7a14 TDn7a28 TDn7a29 1e-9
Ln7a15 TDn7a30 TDn7a31 1e-9
Ln7a16 TDn7a32 TDn7a33 1e-9
Ln8a1 TDn8a2 TDn8a3 1e-9
Ln8a2 TDn8a4 TDn8a5 1e-9
Ln8a3 TDn8a6 TDn8a7 1e-9
Ln8a4 TDn8a8 TDn8a9 1e-9
Ln8a5 TDn8a10 TDn8a11 1e-9
Ln8a6 TDn8a12 TDn8a13 1e-9
Ln8a7 TDn8a14 TDn8a15 1e-9
Ln8a8 TDn8a16 TDn8a17 1e-9
Ln8a9 TDn8a18 TDn8a19 1e-9
Ln8a10 TDn8a20 TDn8a21 1e-9
Ln8a11 TDn8a22 TDn8a23 1e-9
Ln8a12 TDn8a24 TDn8a25 1e-9
Ln8a13 TDn8a26 TDn8a27 1e-9
Ln8a14 TDn8a28 TDn8a29 1e-9
Ln8a15 TDn8a30 TDn8a31 1e-9
Ln8a16 TDn8a32 TDn8a33 1e-9
Ln9a1 TDn9a2 TDn9a3 1e-9
Ln9a2 TDn9a4 TDn9a5 1e-9
Ln9a3 TDn9a6 TDn9a7 1e-9
Ln9a4 TDn9a8 TDn9a9 1e-9
Ln9a5 TDn9a10 TDn9a11 1e-9
Ln9a6 TDn9a12 TDn9a13 1e-9
Ln9a7 TDn9a14 TDn9a15 1e-9
Ln9a8 TDn9a16 TDn9a17 1e-9
Ln9a9 TDn9a18 TDn9a19 1e-9
Ln9a10 TDn9a20 TDn9a21 1e-9
Ln9a11 TDn9a22 TDn9a23 1e-9
Ln9a12 TDn9a24 TDn9a25 1e-9
Ln9a13 TDn9a26 TDn9a27 1e-9
Ln9a14 TDn9a28 TDn9a29 1e-9
Ln9a15 TDn9a30 TDn9a31 1e-9
Ln9a16 TDn9a32 TDn9a33 1e-9
Ln10a1 TDn10a2 TDn10a3 1e-9
Ln10a2 TDn10a4 TDn10a5 1e-9
Ln10a3 TDn10a6 TDn10a7 1e-9
Ln10a4 TDn10a8 TDn10a9 1e-9
Ln10a5 TDn10a10 TDn10a11 1e-9
Ln10a6 TDn10a12 TDn10a13 1e-9
Ln10a7 TDn10a14 TDn10a15 1e-9
Ln10a8 TDn10a16 TDn10a17 1e-9
Ln10a9 TDn10a18 TDn10a19 1e-9
Ln10a10 TDn10a20 TDn10a21 1e-9
Ln10a11 TDn10a22 TDn10a23 1e-9
Ln10a12 TDn10a24 TDn10a25 1e-9
Ln10a13 TDn10a26 TDn10a27 1e-9
Ln10a14 TDn10a28 TDn10a29 1e-9
Ln10a15 TDn10a30 TDn10a31 1e-9
Ln10a16 TDn10a32 TDn10a33 1e-9
Ln11a1 TDn11a2 TDn11a3 1e-9
Ln11a2 TDn11a4 TDn11a5 1e-9
Ln11a3 TDn11a6 TDn11a7 1e-9
Ln11a4 TDn11a8 TDn11a9 1e-9
Ln11a5 TDn11a10 TDn11a11 1e-9
Ln11a6 TDn11a12 TDn11a13 1e-9
Ln11a7 TDn11a14 TDn11a15 1e-9
Ln11a8 TDn11a16 TDn11a17 1e-9
Ln11a9 TDn11a18 TDn11a19 1e-9
Ln11a10 TDn11a20 TDn11a21 1e-9
Ln11a11 TDn11a22 TDn11a23 1e-9
Ln11a12 TDn11a24 TDn11a25 1e-9
Ln11a13 TDn11a26 TDn11a27 1e-9
Ln11a14 TDn11a28 TDn11a29 1e-9
Ln11a15 TDn11a30 TDn11a31 1e-9
Ln11a16 TDn11a32 TDn11a33 1e-9
Ln12a1 TDn12a2 TDn12a3 1e-9
Ln12a2 TDn12a4 TDn12a5 1e-9
Ln12a3 TDn12a6 TDn12a7 1e-9
Ln12a4 TDn12a8 TDn12a9 1e-9
Ln12a5 TDn12a10 TDn12a11 1e-9
Ln12a6 TDn12a12 TDn12a13 1e-9
Ln12a7 TDn12a14 TDn12a15 1e-9
Ln12a8 TDn12a16 TDn12a17 1e-9
Ln12a9 TDn12a18 TDn12a19 1e-9
Ln12a10 TDn12a20 TDn12a21 1e-9
Ln12a11 TDn12a22 TDn12a23 1e-9
Ln12a12 TDn12a24 TDn12a25 1e-9
Ln12a13 TDn12a26 TDn12a27 1e-9
Ln12a14 TDn12a28 TDn12a29 1e-9
Ln12a15 TDn12a30 TDn12a31 1e-9
Ln12a16 TDn12a32 TDn12a33 1e-9
Lnva1 TDnva2 TDnva3 1e-9
Lnva2 TDnva4 TDnva5 1e-9
Lnva3 TDnva6 TDnva7 1e-9
Lnva4 TDnva8 TDnva9 1e-9
Lnva5 TDnva10 TDnva11 1e-9
Lnva6 TDnva12 TDnva13 1e-9
Lnva7 TDnva14 TDnva15 1e-9
Lnva8 TDnva16 TDnva17 1e-9
Lnva9 TDnva18 TDnva19 1e-9
Lnva10 TDnva20 TDnva21 1e-9
Lnva11 TDnva22 TDnva23 1e-9
Lnva12 TDnva24 TDnva25 1e-9
Lnva13 TDnva26 TDnva27 1e-9
Lnva14 TDnva28 TDnva29 1e-9
Lnva15 TDnva30 TDnva31 1e-9
Lnva16 TDnva32 TDnva33 1e-9
Kngan1a1 Lnga1 Ln1a1 0.8
Kngan1a2 Lnga2 Ln1a2 0.8
Kngan1a3 Lnga3 Ln1a3 0.8
Kngan1a4 Lnga4 Ln1a4 0.8
Kngan1a5 Lnga5 Ln1a5 0.8
Kngan1a6 Lnga6 Ln1a6 0.8
Kngan1a7 Lnga7 Ln1a7 0.8
Kngan1a8 Lnga8 Ln1a8 0.8
Kngan1a9 Lnga9 Ln1a9 0.8
Kngan1a10 Lnga10 Ln1a10 0.8
Kngan1a11 Lnga11 Ln1a11 0.8
Kngan1a12 Lnga12 Ln1a12 0.8
Kngan1a13 Lnga13 Ln1a13 0.8
Kngan1a14 Lnga14 Ln1a14 0.8
Kngan1a15 Lnga15 Ln1a15 0.8
Kngan1a16 Lnga16 Ln1a16 0.8
Kngan2a1 Lnga1 Ln2a1 0.7
Kngan2a2 Lnga2 Ln2a2 0.7
Kngan2a3 Lnga3 Ln2a3 0.7
Kngan2a4 Lnga4 Ln2a4 0.7
Kngan2a5 Lnga5 Ln2a5 0.7
Kngan2a6 Lnga6 Ln2a6 0.7
Kngan2a7 Lnga7 Ln2a7 0.7
Kngan2a8 Lnga8 Ln2a8 0.7
Kngan2a9 Lnga9 Ln2a9 0.7
Kngan2a10 Lnga10 Ln2a10 0.7
Kngan2a11 Lnga11 Ln2a11 0.7
Kngan2a12 Lnga12 Ln2a12 0.7
Kngan2a13 Lnga13 Ln2a13 0.7
Kngan2a14 Lnga14 Ln2a14 0.7
Kngan2a15 Lnga15 Ln2a15 0.7
Kngan2a16 Lnga16 Ln2a16 0.7
Kngan3a1 Lnga1 Ln3a1 0.7
Kngan3a2 Lnga2 Ln3a2 0.7
Kngan3a3 Lnga3 Ln3a3 0.7
Kngan3a4 Lnga4 Ln3a4 0.7
Kngan3a5 Lnga5 Ln3a5 0.7
Kngan3a6 Lnga6 Ln3a6 0.7
Kngan3a7 Lnga7 Ln3a7 0.7
Kngan3a8 Lnga8 Ln3a8 0.7
Kngan3a9 Lnga9 Ln3a9 0.7
Kngan3a10 Lnga10 Ln3a10 0.7
Kngan3a11 Lnga11 Ln3a11 0.7
Kngan3a12 Lnga12 Ln3a12 0.7
Kngan3a13 Lnga13 Ln3a13 0.7
Kngan3a14 Lnga14 Ln3a14 0.7
Kngan3a15 Lnga15 Ln3a15 0.7
Kngan3a16 Lnga16 Ln3a16 0.7
Kngan4a1 Lnga1 Ln4a1 0.6
Kngan4a2 Lnga2 Ln4a2 0.6
Kngan4a3 Lnga3 Ln4a3 0.6
Kngan4a4 Lnga4 Ln4a4 0.6
Kngan4a5 Lnga5 Ln4a5 0.6
Kngan4a6 Lnga6 Ln4a6 0.6
Kngan4a7 Lnga7 Ln4a7 0.6
Kngan4a8 Lnga8 Ln4a8 0.6
Kngan4a9 Lnga9 Ln4a9 0.6
Kngan4a10 Lnga10 Ln4a10 0.6
Kngan4a11 Lnga11 Ln4a11 0.6
Kngan4a12 Lnga12 Ln4a12 0.6
Kngan4a13 Lnga13 Ln4a13 0.6
Kngan4a14 Lnga14 Ln4a14 0.6
Kngan4a15 Lnga15 Ln4a15 0.6
Kngan4a16 Lnga16 Ln4a16 0.6
Kngan5a1 Lnga1 Ln5a1 0.6
Kngan5a2 Lnga2 Ln5a2 0.6
Kngan5a3 Lnga3 Ln5a3 0.6
Kngan5a4 Lnga4 Ln5a4 0.6
Kngan5a5 Lnga5 Ln5a5 0.6
Kngan5a6 Lnga6 Ln5a6 0.6
Kngan5a7 Lnga7 Ln5a7 0.6
Kngan5a8 Lnga8 Ln5a8 0.6
Kngan5a9 Lnga9 Ln5a9 0.6
Kngan5a10 Lnga10 Ln5a10 0.6
Kngan5a11 Lnga11 Ln5a11 0.6
Kngan5a12 Lnga12 Ln5a12 0.6
Kngan5a13 Lnga13 Ln5a13 0.6
Kngan5a14 Lnga14 Ln5a14 0.6
Kngan5a15 Lnga15 Ln5a15 0.6
Kngan5a16 Lnga16 Ln5a16 0.6
Kngan6a1 Lnga1 Ln6a1 0.6
Kngan6a2 Lnga2 Ln6a2 0.6
Kngan6a3 Lnga3 Ln6a3 0.6
Kngan6a4 Lnga4 Ln6a4 0.6
Kngan6a5 Lnga5 Ln6a5 0.6
Kngan6a6 Lnga6 Ln6a6 0.6
Kngan6a7 Lnga7 Ln6a7 0.6
Kngan6a8 Lnga8 Ln6a8 0.6
Kngan6a9 Lnga9 Ln6a9 0.6
Kngan6a10 Lnga10 Ln6a10 0.6
Kngan6a11 Lnga11 Ln6a11 0.6
Kngan6a12 Lnga12 Ln6a12 0.6
Kngan6a13 Lnga13 Ln6a13 0.6
Kngan6a14 Lnga14 Ln6a14 0.6
Kngan6a15 Lnga15 Ln6a15 0.6
Kngan6a16 Lnga16 Ln6a16 0.6
Kngan7a1 Lnga1 Ln7a1 0.6
Kngan7a2 Lnga2 Ln7a2 0.6
Kngan7a3 Lnga3 Ln7a3 0.6
Kngan7a4 Lnga4 Ln7a4 0.6
Kngan7a5 Lnga5 Ln7a5 0.6
Kngan7a6 Lnga6 Ln7a6 0.6
Kngan7a7 Lnga7 Ln7a7 0.6
Kngan7a8 Lnga8 Ln7a8 0.6
Kngan7a9 Lnga9 Ln7a9 0.6
Kngan7a10 Lnga10 Ln7a10 0.6
Kngan7a11 Lnga11 Ln7a11 0.6
Kngan7a12 Lnga12 Ln7a12 0.6
Kngan7a13 Lnga13 Ln7a13 0.6
Kngan7a14 Lnga14 Ln7a14 0.6
Kngan7a15 Lnga15 Ln7a15 0.6
Kngan7a16 Lnga16 Ln7a16 0.6
Kngan8a1 Lnga1 Ln8a1 0.6
Kngan8a2 Lnga2 Ln8a2 0.6
Kngan8a3 Lnga3 Ln8a3 0.6
Kngan8a4 Lnga4 Ln8a4 0.6
Kngan8a5 Lnga5 Ln8a5 0.6
Kngan8a6 Lnga6 Ln8a6 0.6
Kngan8a7 Lnga7 Ln8a7 0.6
Kngan8a8 Lnga8 Ln8a8 0.6
Kngan8a9 Lnga9 Ln8a9 0.6
Kngan8a10 Lnga10 Ln8a10 0.6
Kngan8a11 Lnga11 Ln8a11 0.6
Kngan8a12 Lnga12 Ln8a12 0.6
Kngan8a13 Lnga13 Ln8a13 0.6
Kngan8a14 Lnga14 Ln8a14 0.6
Kngan8a15 Lnga15 Ln8a15 0.6
Kngan8a16 Lnga16 Ln8a16 0.6
Kngan9a1 Lnga1 Ln9a1 0.5
Kngan9a2 Lnga2 Ln9a2 0.5
Kngan9a3 Lnga3 Ln9a3 0.5
Kngan9a4 Lnga4 Ln9a4 0.5
Kngan9a5 Lnga5 Ln9a5 0.5
Kngan9a6 Lnga6 Ln9a6 0.5
Kngan9a7 Lnga7 Ln9a7 0.5
Kngan9a8 Lnga8 Ln9a8 0.5
Kngan9a9 Lnga9 Ln9a9 0.5
Kngan9a10 Lnga10 Ln9a10 0.5
Kngan9a11 Lnga11 Ln9a11 0.5
Kngan9a12 Lnga12 Ln9a12 0.5
Kngan9a13 Lnga13 Ln9a13 0.5
Kngan9a14 Lnga14 Ln9a14 0.5
Kngan9a15 Lnga15 Ln9a15 0.5
Kngan9a16 Lnga16 Ln9a16 0.5
Kngan10a1 Lnga1 Ln10a1 0.5
Kngan10a2 Lnga2 Ln10a2 0.5
Kngan10a3 Lnga3 Ln10a3 0.5
Kngan10a4 Lnga4 Ln10a4 0.5
Kngan10a5 Lnga5 Ln10a5 0.5
Kngan10a6 Lnga6 Ln10a6 0.5
Kngan10a7 Lnga7 Ln10a7 0.5
Kngan10a8 Lnga8 Ln10a8 0.5
Kngan10a9 Lnga9 Ln10a9 0.5
Kngan10a10 Lnga10 Ln10a10 0.5
Kngan10a11 Lnga11 Ln10a11 0.5
Kngan10a12 Lnga12 Ln10a12 0.5
Kngan10a13 Lnga13 Ln10a13 0.5
Kngan10a14 Lnga14 Ln10a14 0.5
Kngan10a15 Lnga15 Ln10a15 0.5
Kngan10a16 Lnga16 Ln10a16 0.5
Kngan11a1 Lnga1 Ln11a1 0.5
Kngan11a2 Lnga2 Ln11a2 0.5
Kngan11a3 Lnga3 Ln11a3 0.5
Kngan11a4 Lnga4 Ln11a4 0.5
Kngan11a5 Lnga5 Ln11a5 0.5
Kngan11a6 Lnga6 Ln11a6 0.5
Kngan11a7 Lnga7 Ln11a7 0.5
Kngan11a8 Lnga8 Ln11a8 0.5
Kngan11a9 Lnga9 Ln11a9 0.5
Kngan11a10 Lnga10 Ln11a10 0.5
Kngan11a11 Lnga11 Ln11a11 0.5
Kngan11a12 Lnga12 Ln11a12 0.5
Kngan11a13 Lnga13 Ln11a13 0.5
Kngan11a14 Lnga14 Ln11a14 0.5
Kngan11a15 Lnga15 Ln11a15 0.5
Kngan11a16 Lnga16 Ln11a16 0.5
Kngan12a1 Lnga1 Ln12a1 0.5
Kngan12a2 Lnga2 Ln12a2 0.5
Kngan12a3 Lnga3 Ln12a3 0.5
Kngan12a4 Lnga4 Ln12a4 0.5
Kngan12a5 Lnga5 Ln12a5 0.5
Kngan12a6 Lnga6 Ln12a6 0.5
Kngan12a7 Lnga7 Ln12a7 0.5
Kngan12a8 Lnga8 Ln12a8 0.5
Kngan12a9 Lnga9 Ln12a9 0.5
Kngan12a10 Lnga10 Ln12a10 0.5
Kngan12a11 Lnga11 Ln12a11 0.5
Kngan12a12 Lnga12 Ln12a12 0.5
Kngan12a13 Lnga13 Ln12a13 0.5
Kngan12a14 Lnga14 Ln12a14 0.5
Kngan12a15 Lnga15 Ln12a15 0.5
Kngan12a16 Lnga16 Ln12a16 0.5
Knganva1 Lnga1 Lnva1 0.5
Knganva2 Lnga2 Lnva2 0.5
Knganva3 Lnga3 Lnva3 0.5
Knganva4 Lnga4 Lnva4 0.5
Knganva5 Lnga5 Lnva5 0.5
Knganva6 Lnga6 Lnva6 0.5
Knganva7 Lnga7 Lnva7 0.5
Knganva8 Lnga8 Lnva8 0.5
Knganva9 Lnga9 Lnva9 0.5
Knganva10 Lnga10 Lnva10 0.5
Knganva11 Lnga11 Lnva11 0.5
Knganva12 Lnga12 Lnva12 0.5
Knganva13 Lnga13 Lnva13 0.5
Knganva14 Lnga14 Lnva14 0.5
Knganva15 Lnga15 Lnva15 0.5
Knganva16 Lnga16 Lnva16 0.5
Kn1an2a1 Ln1a1 Ln2a1 0.8
Kn1an2a2 Ln1a2 Ln2a2 0.8
Kn1an2a3 Ln1a3 Ln2a3 0.8
Kn1an2a4 Ln1a4 Ln2a4 0.8
Kn1an2a5 Ln1a5 Ln2a5 0.8
Kn1an2a6 Ln1a6 Ln2a6 0.8
Kn1an2a7 Ln1a7 Ln2a7 0.8
Kn1an2a8 Ln1a8 Ln2a8 0.8
Kn1an2a9 Ln1a9 Ln2a9 0.8
Kn1an2a10 Ln1a10 Ln2a10 0.8
Kn1an2a11 Ln1a11 Ln2a11 0.8
Kn1an2a12 Ln1a12 Ln2a12 0.8
Kn1an2a13 Ln1a13 Ln2a13 0.8
Kn1an2a14 Ln1a14 Ln2a14 0.8
Kn1an2a15 Ln1a15 Ln2a15 0.8
Kn1an2a16 Ln1a16 Ln2a16 0.8
Kn1an3a1 Ln1a1 Ln3a1 0.7
Kn1an3a2 Ln1a2 Ln3a2 0.7
Kn1an3a3 Ln1a3 Ln3a3 0.7
Kn1an3a4 Ln1a4 Ln3a4 0.7
Kn1an3a5 Ln1a5 Ln3a5 0.7
Kn1an3a6 Ln1a6 Ln3a6 0.7
Kn1an3a7 Ln1a7 Ln3a7 0.7
Kn1an3a8 Ln1a8 Ln3a8 0.7
Kn1an3a9 Ln1a9 Ln3a9 0.7
Kn1an3a10 Ln1a10 Ln3a10 0.7
Kn1an3a11 Ln1a11 Ln3a11 0.7
Kn1an3a12 Ln1a12 Ln3a12 0.7
Kn1an3a13 Ln1a13 Ln3a13 0.7
Kn1an3a14 Ln1a14 Ln3a14 0.7
Kn1an3a15 Ln1a15 Ln3a15 0.7
Kn1an3a16 Ln1a16 Ln3a16 0.7
Kn1an4a1 Ln1a1 Ln4a1 0.7
Kn1an4a2 Ln1a2 Ln4a2 0.7
Kn1an4a3 Ln1a3 Ln4a3 0.7
Kn1an4a4 Ln1a4 Ln4a4 0.7
Kn1an4a5 Ln1a5 Ln4a5 0.7
Kn1an4a6 Ln1a6 Ln4a6 0.7
Kn1an4a7 Ln1a7 Ln4a7 0.7
Kn1an4a8 Ln1a8 Ln4a8 0.7
Kn1an4a9 Ln1a9 Ln4a9 0.7
Kn1an4a10 Ln1a10 Ln4a10 0.7
Kn1an4a11 Ln1a11 Ln4a11 0.7
Kn1an4a12 Ln1a12 Ln4a12 0.7
Kn1an4a13 Ln1a13 Ln4a13 0.7
Kn1an4a14 Ln1a14 Ln4a14 0.7
Kn1an4a15 Ln1a15 Ln4a15 0.7
Kn1an4a16 Ln1a16 Ln4a16 0.7
Kn1an5a1 Ln1a1 Ln5a1 0.6
Kn1an5a2 Ln1a2 Ln5a2 0.6
Kn1an5a3 Ln1a3 Ln5a3 0.6
Kn1an5a4 Ln1a4 Ln5a4 0.6
Kn1an5a5 Ln1a5 Ln5a5 0.6
Kn1an5a6 Ln1a6 Ln5a6 0.6
Kn1an5a7 Ln1a7 Ln5a7 0.6
Kn1an5a8 Ln1a8 Ln5a8 0.6
Kn1an5a9 Ln1a9 Ln5a9 0.6
Kn1an5a10 Ln1a10 Ln5a10 0.6
Kn1an5a11 Ln1a11 Ln5a11 0.6
Kn1an5a12 Ln1a12 Ln5a12 0.6
Kn1an5a13 Ln1a13 Ln5a13 0.6
Kn1an5a14 Ln1a14 Ln5a14 0.6
Kn1an5a15 Ln1a15 Ln5a15 0.6
Kn1an5a16 Ln1a16 Ln5a16 0.6
Kn1an6a1 Ln1a1 Ln6a1 0.6
Kn1an6a2 Ln1a2 Ln6a2 0.6
Kn1an6a3 Ln1a3 Ln6a3 0.6
Kn1an6a4 Ln1a4 Ln6a4 0.6
Kn1an6a5 Ln1a5 Ln6a5 0.6
Kn1an6a6 Ln1a6 Ln6a6 0.6
Kn1an6a7 Ln1a7 Ln6a7 0.6
Kn1an6a8 Ln1a8 Ln6a8 0.6
Kn1an6a9 Ln1a9 Ln6a9 0.6
Kn1an6a10 Ln1a10 Ln6a10 0.6
Kn1an6a11 Ln1a11 Ln6a11 0.6
Kn1an6a12 Ln1a12 Ln6a12 0.6
Kn1an6a13 Ln1a13 Ln6a13 0.6
Kn1an6a14 Ln1a14 Ln6a14 0.6
Kn1an6a15 Ln1a15 Ln6a15 0.6
Kn1an6a16 Ln1a16 Ln6a16 0.6
Kn1an7a1 Ln1a1 Ln7a1 0.6
Kn1an7a2 Ln1a2 Ln7a2 0.6
Kn1an7a3 Ln1a3 Ln7a3 0.6
Kn1an7a4 Ln1a4 Ln7a4 0.6
Kn1an7a5 Ln1a5 Ln7a5 0.6
Kn1an7a6 Ln1a6 Ln7a6 0.6
Kn1an7a7 Ln1a7 Ln7a7 0.6
Kn1an7a8 Ln1a8 Ln7a8 0.6
Kn1an7a9 Ln1a9 Ln7a9 0.6
Kn1an7a10 Ln1a10 Ln7a10 0.6
Kn1an7a11 Ln1a11 Ln7a11 0.6
Kn1an7a12 Ln1a12 Ln7a12 0.6
Kn1an7a13 Ln1a13 Ln7a13 0.6
Kn1an7a14 Ln1a14 Ln7a14 0.6
Kn1an7a15 Ln1a15 Ln7a15 0.6
Kn1an7a16 Ln1a16 Ln7a16 0.6
Kn1an8a1 Ln1a1 Ln8a1 0.6
Kn1an8a2 Ln1a2 Ln8a2 0.6
Kn1an8a3 Ln1a3 Ln8a3 0.6
Kn1an8a4 Ln1a4 Ln8a4 0.6
Kn1an8a5 Ln1a5 Ln8a5 0.6
Kn1an8a6 Ln1a6 Ln8a6 0.6
Kn1an8a7 Ln1a7 Ln8a7 0.6
Kn1an8a8 Ln1a8 Ln8a8 0.6
Kn1an8a9 Ln1a9 Ln8a9 0.6
Kn1an8a10 Ln1a10 Ln8a10 0.6
Kn1an8a11 Ln1a11 Ln8a11 0.6
Kn1an8a12 Ln1a12 Ln8a12 0.6
Kn1an8a13 Ln1a13 Ln8a13 0.6
Kn1an8a14 Ln1a14 Ln8a14 0.6
Kn1an8a15 Ln1a15 Ln8a15 0.6
Kn1an8a16 Ln1a16 Ln8a16 0.6
Kn1an9a1 Ln1a1 Ln9a1 0.6
Kn1an9a2 Ln1a2 Ln9a2 0.6
Kn1an9a3 Ln1a3 Ln9a3 0.6
Kn1an9a4 Ln1a4 Ln9a4 0.6
Kn1an9a5 Ln1a5 Ln9a5 0.6
Kn1an9a6 Ln1a6 Ln9a6 0.6
Kn1an9a7 Ln1a7 Ln9a7 0.6
Kn1an9a8 Ln1a8 Ln9a8 0.6
Kn1an9a9 Ln1a9 Ln9a9 0.6
Kn1an9a10 Ln1a10 Ln9a10 0.6
Kn1an9a11 Ln1a11 Ln9a11 0.6
Kn1an9a12 Ln1a12 Ln9a12 0.6
Kn1an9a13 Ln1a13 Ln9a13 0.6
Kn1an9a14 Ln1a14 Ln9a14 0.6
Kn1an9a15 Ln1a15 Ln9a15 0.6
Kn1an9a16 Ln1a16 Ln9a16 0.6
Kn1an10a1 Ln1a1 Ln10a1 0.5
Kn1an10a2 Ln1a2 Ln10a2 0.5
Kn1an10a3 Ln1a3 Ln10a3 0.5
Kn1an10a4 Ln1a4 Ln10a4 0.5
Kn1an10a5 Ln1a5 Ln10a5 0.5
Kn1an10a6 Ln1a6 Ln10a6 0.5
Kn1an10a7 Ln1a7 Ln10a7 0.5
Kn1an10a8 Ln1a8 Ln10a8 0.5
Kn1an10a9 Ln1a9 Ln10a9 0.5
Kn1an10a10 Ln1a10 Ln10a10 0.5
Kn1an10a11 Ln1a11 Ln10a11 0.5
Kn1an10a12 Ln1a12 Ln10a12 0.5
Kn1an10a13 Ln1a13 Ln10a13 0.5
Kn1an10a14 Ln1a14 Ln10a14 0.5
Kn1an10a15 Ln1a15 Ln10a15 0.5
Kn1an10a16 Ln1a16 Ln10a16 0.5
Kn1an11a1 Ln1a1 Ln11a1 0.5
Kn1an11a2 Ln1a2 Ln11a2 0.5
Kn1an11a3 Ln1a3 Ln11a3 0.5
Kn1an11a4 Ln1a4 Ln11a4 0.5
Kn1an11a5 Ln1a5 Ln11a5 0.5
Kn1an11a6 Ln1a6 Ln11a6 0.5
Kn1an11a7 Ln1a7 Ln11a7 0.5
Kn1an11a8 Ln1a8 Ln11a8 0.5
Kn1an11a9 Ln1a9 Ln11a9 0.5
Kn1an11a10 Ln1a10 Ln11a10 0.5
Kn1an11a11 Ln1a11 Ln11a11 0.5
Kn1an11a12 Ln1a12 Ln11a12 0.5
Kn1an11a13 Ln1a13 Ln11a13 0.5
Kn1an11a14 Ln1a14 Ln11a14 0.5
Kn1an11a15 Ln1a15 Ln11a15 0.5
Kn1an11a16 Ln1a16 Ln11a16 0.5
Kn1an12a1 Ln1a1 Ln12a1 0.5
Kn1an12a2 Ln1a2 Ln12a2 0.5
Kn1an12a3 Ln1a3 Ln12a3 0.5
Kn1an12a4 Ln1a4 Ln12a4 0.5
Kn1an12a5 Ln1a5 Ln12a5 0.5
Kn1an12a6 Ln1a6 Ln12a6 0.5
Kn1an12a7 Ln1a7 Ln12a7 0.5
Kn1an12a8 Ln1a8 Ln12a8 0.5
Kn1an12a9 Ln1a9 Ln12a9 0.5
Kn1an12a10 Ln1a10 Ln12a10 0.5
Kn1an12a11 Ln1a11 Ln12a11 0.5
Kn1an12a12 Ln1a12 Ln12a12 0.5
Kn1an12a13 Ln1a13 Ln12a13 0.5
Kn1an12a14 Ln1a14 Ln12a14 0.5
Kn1an12a15 Ln1a15 Ln12a15 0.5
Kn1an12a16 Ln1a16 Ln12a16 0.5
Kn1anva1 Ln1a1 Lnva1 0.5
Kn1anva2 Ln1a2 Lnva2 0.5
Kn1anva3 Ln1a3 Lnva3 0.5
Kn1anva4 Ln1a4 Lnva4 0.5
Kn1anva5 Ln1a5 Lnva5 0.5
Kn1anva6 Ln1a6 Lnva6 0.5
Kn1anva7 Ln1a7 Lnva7 0.5
Kn1anva8 Ln1a8 Lnva8 0.5
Kn1anva9 Ln1a9 Lnva9 0.5
Kn1anva10 Ln1a10 Lnva10 0.5
Kn1anva11 Ln1a11 Lnva11 0.5
Kn1anva12 Ln1a12 Lnva12 0.5
Kn1anva13 Ln1a13 Lnva13 0.5
Kn1anva14 Ln1a14 Lnva14 0.5
Kn1anva15 Ln1a15 Lnva15 0.5
Kn1anva16 Ln1a16 Lnva16 0.5
Kn2an3a1 Ln2a1 Ln3a1 0.8
Kn2an3a2 Ln2a2 Ln3a2 0.8
Kn2an3a3 Ln2a3 Ln3a3 0.8
Kn2an3a4 Ln2a4 Ln3a4 0.8
Kn2an3a5 Ln2a5 Ln3a5 0.8
Kn2an3a6 Ln2a6 Ln3a6 0.8
Kn2an3a7 Ln2a7 Ln3a7 0.8
Kn2an3a8 Ln2a8 Ln3a8 0.8
Kn2an3a9 Ln2a9 Ln3a9 0.8
Kn2an3a10 Ln2a10 Ln3a10 0.8
Kn2an3a11 Ln2a11 Ln3a11 0.8
Kn2an3a12 Ln2a12 Ln3a12 0.8
Kn2an3a13 Ln2a13 Ln3a13 0.8
Kn2an3a14 Ln2a14 Ln3a14 0.8
Kn2an3a15 Ln2a15 Ln3a15 0.8
Kn2an3a16 Ln2a16 Ln3a16 0.8
Kn2an4a1 Ln2a1 Ln4a1 0.7
Kn2an4a2 Ln2a2 Ln4a2 0.7
Kn2an4a3 Ln2a3 Ln4a3 0.7
Kn2an4a4 Ln2a4 Ln4a4 0.7
Kn2an4a5 Ln2a5 Ln4a5 0.7
Kn2an4a6 Ln2a6 Ln4a6 0.7
Kn2an4a7 Ln2a7 Ln4a7 0.7
Kn2an4a8 Ln2a8 Ln4a8 0.7
Kn2an4a9 Ln2a9 Ln4a9 0.7
Kn2an4a10 Ln2a10 Ln4a10 0.7
Kn2an4a11 Ln2a11 Ln4a11 0.7
Kn2an4a12 Ln2a12 Ln4a12 0.7
Kn2an4a13 Ln2a13 Ln4a13 0.7
Kn2an4a14 Ln2a14 Ln4a14 0.7
Kn2an4a15 Ln2a15 Ln4a15 0.7
Kn2an4a16 Ln2a16 Ln4a16 0.7
Kn2an5a1 Ln2a1 Ln5a1 0.7
Kn2an5a2 Ln2a2 Ln5a2 0.7
Kn2an5a3 Ln2a3 Ln5a3 0.7
Kn2an5a4 Ln2a4 Ln5a4 0.7
Kn2an5a5 Ln2a5 Ln5a5 0.7
Kn2an5a6 Ln2a6 Ln5a6 0.7
Kn2an5a7 Ln2a7 Ln5a7 0.7
Kn2an5a8 Ln2a8 Ln5a8 0.7
Kn2an5a9 Ln2a9 Ln5a9 0.7
Kn2an5a10 Ln2a10 Ln5a10 0.7
Kn2an5a11 Ln2a11 Ln5a11 0.7
Kn2an5a12 Ln2a12 Ln5a12 0.7
Kn2an5a13 Ln2a13 Ln5a13 0.7
Kn2an5a14 Ln2a14 Ln5a14 0.7
Kn2an5a15 Ln2a15 Ln5a15 0.7
Kn2an5a16 Ln2a16 Ln5a16 0.7
Kn2an6a1 Ln2a1 Ln6a1 0.6
Kn2an6a2 Ln2a2 Ln6a2 0.6
Kn2an6a3 Ln2a3 Ln6a3 0.6
Kn2an6a4 Ln2a4 Ln6a4 0.6
Kn2an6a5 Ln2a5 Ln6a5 0.6
Kn2an6a6 Ln2a6 Ln6a6 0.6
Kn2an6a7 Ln2a7 Ln6a7 0.6
Kn2an6a8 Ln2a8 Ln6a8 0.6
Kn2an6a9 Ln2a9 Ln6a9 0.6
Kn2an6a10 Ln2a10 Ln6a10 0.6
Kn2an6a11 Ln2a11 Ln6a11 0.6
Kn2an6a12 Ln2a12 Ln6a12 0.6
Kn2an6a13 Ln2a13 Ln6a13 0.6
Kn2an6a14 Ln2a14 Ln6a14 0.6
Kn2an6a15 Ln2a15 Ln6a15 0.6
Kn2an6a16 Ln2a16 Ln6a16 0.6
Kn2an7a1 Ln2a1 Ln7a1 0.6
Kn2an7a2 Ln2a2 Ln7a2 0.6
Kn2an7a3 Ln2a3 Ln7a3 0.6
Kn2an7a4 Ln2a4 Ln7a4 0.6
Kn2an7a5 Ln2a5 Ln7a5 0.6
Kn2an7a6 Ln2a6 Ln7a6 0.6
Kn2an7a7 Ln2a7 Ln7a7 0.6
Kn2an7a8 Ln2a8 Ln7a8 0.6
Kn2an7a9 Ln2a9 Ln7a9 0.6
Kn2an7a10 Ln2a10 Ln7a10 0.6
Kn2an7a11 Ln2a11 Ln7a11 0.6
Kn2an7a12 Ln2a12 Ln7a12 0.6
Kn2an7a13 Ln2a13 Ln7a13 0.6
Kn2an7a14 Ln2a14 Ln7a14 0.6
Kn2an7a15 Ln2a15 Ln7a15 0.6
Kn2an7a16 Ln2a16 Ln7a16 0.6
Kn2an8a1 Ln2a1 Ln8a1 0.6
Kn2an8a2 Ln2a2 Ln8a2 0.6
Kn2an8a3 Ln2a3 Ln8a3 0.6
Kn2an8a4 Ln2a4 Ln8a4 0.6
Kn2an8a5 Ln2a5 Ln8a5 0.6
Kn2an8a6 Ln2a6 Ln8a6 0.6
Kn2an8a7 Ln2a7 Ln8a7 0.6
Kn2an8a8 Ln2a8 Ln8a8 0.6
Kn2an8a9 Ln2a9 Ln8a9 0.6
Kn2an8a10 Ln2a10 Ln8a10 0.6
Kn2an8a11 Ln2a11 Ln8a11 0.6
Kn2an8a12 Ln2a12 Ln8a12 0.6
Kn2an8a13 Ln2a13 Ln8a13 0.6
Kn2an8a14 Ln2a14 Ln8a14 0.6
Kn2an8a15 Ln2a15 Ln8a15 0.6
Kn2an8a16 Ln2a16 Ln8a16 0.6
Kn2an9a1 Ln2a1 Ln9a1 0.6
Kn2an9a2 Ln2a2 Ln9a2 0.6
Kn2an9a3 Ln2a3 Ln9a3 0.6
Kn2an9a4 Ln2a4 Ln9a4 0.6
Kn2an9a5 Ln2a5 Ln9a5 0.6
Kn2an9a6 Ln2a6 Ln9a6 0.6
Kn2an9a7 Ln2a7 Ln9a7 0.6
Kn2an9a8 Ln2a8 Ln9a8 0.6
Kn2an9a9 Ln2a9 Ln9a9 0.6
Kn2an9a10 Ln2a10 Ln9a10 0.6
Kn2an9a11 Ln2a11 Ln9a11 0.6
Kn2an9a12 Ln2a12 Ln9a12 0.6
Kn2an9a13 Ln2a13 Ln9a13 0.6
Kn2an9a14 Ln2a14 Ln9a14 0.6
Kn2an9a15 Ln2a15 Ln9a15 0.6
Kn2an9a16 Ln2a16 Ln9a16 0.6
Kn2an10a1 Ln2a1 Ln10a1 0.6
Kn2an10a2 Ln2a2 Ln10a2 0.6
Kn2an10a3 Ln2a3 Ln10a3 0.6
Kn2an10a4 Ln2a4 Ln10a4 0.6
Kn2an10a5 Ln2a5 Ln10a5 0.6
Kn2an10a6 Ln2a6 Ln10a6 0.6
Kn2an10a7 Ln2a7 Ln10a7 0.6
Kn2an10a8 Ln2a8 Ln10a8 0.6
Kn2an10a9 Ln2a9 Ln10a9 0.6
Kn2an10a10 Ln2a10 Ln10a10 0.6
Kn2an10a11 Ln2a11 Ln10a11 0.6
Kn2an10a12 Ln2a12 Ln10a12 0.6
Kn2an10a13 Ln2a13 Ln10a13 0.6
Kn2an10a14 Ln2a14 Ln10a14 0.6
Kn2an10a15 Ln2a15 Ln10a15 0.6
Kn2an10a16 Ln2a16 Ln10a16 0.6
Kn2an11a1 Ln2a1 Ln11a1 0.5
Kn2an11a2 Ln2a2 Ln11a2 0.5
Kn2an11a3 Ln2a3 Ln11a3 0.5
Kn2an11a4 Ln2a4 Ln11a4 0.5
Kn2an11a5 Ln2a5 Ln11a5 0.5
Kn2an11a6 Ln2a6 Ln11a6 0.5
Kn2an11a7 Ln2a7 Ln11a7 0.5
Kn2an11a8 Ln2a8 Ln11a8 0.5
Kn2an11a9 Ln2a9 Ln11a9 0.5
Kn2an11a10 Ln2a10 Ln11a10 0.5
Kn2an11a11 Ln2a11 Ln11a11 0.5
Kn2an11a12 Ln2a12 Ln11a12 0.5
Kn2an11a13 Ln2a13 Ln11a13 0.5
Kn2an11a14 Ln2a14 Ln11a14 0.5
Kn2an11a15 Ln2a15 Ln11a15 0.5
Kn2an11a16 Ln2a16 Ln11a16 0.5
Kn2an12a1 Ln2a1 Ln12a1 0.5
Kn2an12a2 Ln2a2 Ln12a2 0.5
Kn2an12a3 Ln2a3 Ln12a3 0.5
Kn2an12a4 Ln2a4 Ln12a4 0.5
Kn2an12a5 Ln2a5 Ln12a5 0.5
Kn2an12a6 Ln2a6 Ln12a6 0.5
Kn2an12a7 Ln2a7 Ln12a7 0.5
Kn2an12a8 Ln2a8 Ln12a8 0.5
Kn2an12a9 Ln2a9 Ln12a9 0.5
Kn2an12a10 Ln2a10 Ln12a10 0.5
Kn2an12a11 Ln2a11 Ln12a11 0.5
Kn2an12a12 Ln2a12 Ln12a12 0.5
Kn2an12a13 Ln2a13 Ln12a13 0.5
Kn2an12a14 Ln2a14 Ln12a14 0.5
Kn2an12a15 Ln2a15 Ln12a15 0.5
Kn2an12a16 Ln2a16 Ln12a16 0.5
Kn2anva1 Ln2a1 Lnva1 0.5
Kn2anva2 Ln2a2 Lnva2 0.5
Kn2anva3 Ln2a3 Lnva3 0.5
Kn2anva4 Ln2a4 Lnva4 0.5
Kn2anva5 Ln2a5 Lnva5 0.5
Kn2anva6 Ln2a6 Lnva6 0.5
Kn2anva7 Ln2a7 Lnva7 0.5
Kn2anva8 Ln2a8 Lnva8 0.5
Kn2anva9 Ln2a9 Lnva9 0.5
Kn2anva10 Ln2a10 Lnva10 0.5
Kn2anva11 Ln2a11 Lnva11 0.5
Kn2anva12 Ln2a12 Lnva12 0.5
Kn2anva13 Ln2a13 Lnva13 0.5
Kn2anva14 Ln2a14 Lnva14 0.5
Kn2anva15 Ln2a15 Lnva15 0.5
Kn2anva16 Ln2a16 Lnva16 0.5
Kn3an4a1 Ln3a1 Ln4a1 0.8
Kn3an4a2 Ln3a2 Ln4a2 0.8
Kn3an4a3 Ln3a3 Ln4a3 0.8
Kn3an4a4 Ln3a4 Ln4a4 0.8
Kn3an4a5 Ln3a5 Ln4a5 0.8
Kn3an4a6 Ln3a6 Ln4a6 0.8
Kn3an4a7 Ln3a7 Ln4a7 0.8
Kn3an4a8 Ln3a8 Ln4a8 0.8
Kn3an4a9 Ln3a9 Ln4a9 0.8
Kn3an4a10 Ln3a10 Ln4a10 0.8
Kn3an4a11 Ln3a11 Ln4a11 0.8
Kn3an4a12 Ln3a12 Ln4a12 0.8
Kn3an4a13 Ln3a13 Ln4a13 0.8
Kn3an4a14 Ln3a14 Ln4a14 0.8
Kn3an4a15 Ln3a15 Ln4a15 0.8
Kn3an4a16 Ln3a16 Ln4a16 0.8
Kn3an5a1 Ln3a1 Ln5a1 0.7
Kn3an5a2 Ln3a2 Ln5a2 0.7
Kn3an5a3 Ln3a3 Ln5a3 0.7
Kn3an5a4 Ln3a4 Ln5a4 0.7
Kn3an5a5 Ln3a5 Ln5a5 0.7
Kn3an5a6 Ln3a6 Ln5a6 0.7
Kn3an5a7 Ln3a7 Ln5a7 0.7
Kn3an5a8 Ln3a8 Ln5a8 0.7
Kn3an5a9 Ln3a9 Ln5a9 0.7
Kn3an5a10 Ln3a10 Ln5a10 0.7
Kn3an5a11 Ln3a11 Ln5a11 0.7
Kn3an5a12 Ln3a12 Ln5a12 0.7
Kn3an5a13 Ln3a13 Ln5a13 0.7
Kn3an5a14 Ln3a14 Ln5a14 0.7
Kn3an5a15 Ln3a15 Ln5a15 0.7
Kn3an5a16 Ln3a16 Ln5a16 0.7
Kn3an6a1 Ln3a1 Ln6a1 0.7
Kn3an6a2 Ln3a2 Ln6a2 0.7
Kn3an6a3 Ln3a3 Ln6a3 0.7
Kn3an6a4 Ln3a4 Ln6a4 0.7
Kn3an6a5 Ln3a5 Ln6a5 0.7
Kn3an6a6 Ln3a6 Ln6a6 0.7
Kn3an6a7 Ln3a7 Ln6a7 0.7
Kn3an6a8 Ln3a8 Ln6a8 0.7
Kn3an6a9 Ln3a9 Ln6a9 0.7
Kn3an6a10 Ln3a10 Ln6a10 0.7
Kn3an6a11 Ln3a11 Ln6a11 0.7
Kn3an6a12 Ln3a12 Ln6a12 0.7
Kn3an6a13 Ln3a13 Ln6a13 0.7
Kn3an6a14 Ln3a14 Ln6a14 0.7
Kn3an6a15 Ln3a15 Ln6a15 0.7
Kn3an6a16 Ln3a16 Ln6a16 0.7
Kn3an7a1 Ln3a1 Ln7a1 0.6
Kn3an7a2 Ln3a2 Ln7a2 0.6
Kn3an7a3 Ln3a3 Ln7a3 0.6
Kn3an7a4 Ln3a4 Ln7a4 0.6
Kn3an7a5 Ln3a5 Ln7a5 0.6
Kn3an7a6 Ln3a6 Ln7a6 0.6
Kn3an7a7 Ln3a7 Ln7a7 0.6
Kn3an7a8 Ln3a8 Ln7a8 0.6
Kn3an7a9 Ln3a9 Ln7a9 0.6
Kn3an7a10 Ln3a10 Ln7a10 0.6
Kn3an7a11 Ln3a11 Ln7a11 0.6
Kn3an7a12 Ln3a12 Ln7a12 0.6
Kn3an7a13 Ln3a13 Ln7a13 0.6
Kn3an7a14 Ln3a14 Ln7a14 0.6
Kn3an7a15 Ln3a15 Ln7a15 0.6
Kn3an7a16 Ln3a16 Ln7a16 0.6
Kn3an8a1 Ln3a1 Ln8a1 0.6
Kn3an8a2 Ln3a2 Ln8a2 0.6
Kn3an8a3 Ln3a3 Ln8a3 0.6
Kn3an8a4 Ln3a4 Ln8a4 0.6
Kn3an8a5 Ln3a5 Ln8a5 0.6
Kn3an8a6 Ln3a6 Ln8a6 0.6
Kn3an8a7 Ln3a7 Ln8a7 0.6
Kn3an8a8 Ln3a8 Ln8a8 0.6
Kn3an8a9 Ln3a9 Ln8a9 0.6
Kn3an8a10 Ln3a10 Ln8a10 0.6
Kn3an8a11 Ln3a11 Ln8a11 0.6
Kn3an8a12 Ln3a12 Ln8a12 0.6
Kn3an8a13 Ln3a13 Ln8a13 0.6
Kn3an8a14 Ln3a14 Ln8a14 0.6
Kn3an8a15 Ln3a15 Ln8a15 0.6
Kn3an8a16 Ln3a16 Ln8a16 0.6
Kn3an9a1 Ln3a1 Ln9a1 0.6
Kn3an9a2 Ln3a2 Ln9a2 0.6
Kn3an9a3 Ln3a3 Ln9a3 0.6
Kn3an9a4 Ln3a4 Ln9a4 0.6
Kn3an9a5 Ln3a5 Ln9a5 0.6
Kn3an9a6 Ln3a6 Ln9a6 0.6
Kn3an9a7 Ln3a7 Ln9a7 0.6
Kn3an9a8 Ln3a8 Ln9a8 0.6
Kn3an9a9 Ln3a9 Ln9a9 0.6
Kn3an9a10 Ln3a10 Ln9a10 0.6
Kn3an9a11 Ln3a11 Ln9a11 0.6
Kn3an9a12 Ln3a12 Ln9a12 0.6
Kn3an9a13 Ln3a13 Ln9a13 0.6
Kn3an9a14 Ln3a14 Ln9a14 0.6
Kn3an9a15 Ln3a15 Ln9a15 0.6
Kn3an9a16 Ln3a16 Ln9a16 0.6
Kn3an10a1 Ln3a1 Ln10a1 0.6
Kn3an10a2 Ln3a2 Ln10a2 0.6
Kn3an10a3 Ln3a3 Ln10a3 0.6
Kn3an10a4 Ln3a4 Ln10a4 0.6
Kn3an10a5 Ln3a5 Ln10a5 0.6
Kn3an10a6 Ln3a6 Ln10a6 0.6
Kn3an10a7 Ln3a7 Ln10a7 0.6
Kn3an10a8 Ln3a8 Ln10a8 0.6
Kn3an10a9 Ln3a9 Ln10a9 0.6
Kn3an10a10 Ln3a10 Ln10a10 0.6
Kn3an10a11 Ln3a11 Ln10a11 0.6
Kn3an10a12 Ln3a12 Ln10a12 0.6
Kn3an10a13 Ln3a13 Ln10a13 0.6
Kn3an10a14 Ln3a14 Ln10a14 0.6
Kn3an10a15 Ln3a15 Ln10a15 0.6
Kn3an10a16 Ln3a16 Ln10a16 0.6
Kn3an11a1 Ln3a1 Ln11a1 0.6
Kn3an11a2 Ln3a2 Ln11a2 0.6
Kn3an11a3 Ln3a3 Ln11a3 0.6
Kn3an11a4 Ln3a4 Ln11a4 0.6
Kn3an11a5 Ln3a5 Ln11a5 0.6
Kn3an11a6 Ln3a6 Ln11a6 0.6
Kn3an11a7 Ln3a7 Ln11a7 0.6
Kn3an11a8 Ln3a8 Ln11a8 0.6
Kn3an11a9 Ln3a9 Ln11a9 0.6
Kn3an11a10 Ln3a10 Ln11a10 0.6
Kn3an11a11 Ln3a11 Ln11a11 0.6
Kn3an11a12 Ln3a12 Ln11a12 0.6
Kn3an11a13 Ln3a13 Ln11a13 0.6
Kn3an11a14 Ln3a14 Ln11a14 0.6
Kn3an11a15 Ln3a15 Ln11a15 0.6
Kn3an11a16 Ln3a16 Ln11a16 0.6
Kn3an12a1 Ln3a1 Ln12a1 0.5
Kn3an12a2 Ln3a2 Ln12a2 0.5
Kn3an12a3 Ln3a3 Ln12a3 0.5
Kn3an12a4 Ln3a4 Ln12a4 0.5
Kn3an12a5 Ln3a5 Ln12a5 0.5
Kn3an12a6 Ln3a6 Ln12a6 0.5
Kn3an12a7 Ln3a7 Ln12a7 0.5
Kn3an12a8 Ln3a8 Ln12a8 0.5
Kn3an12a9 Ln3a9 Ln12a9 0.5
Kn3an12a10 Ln3a10 Ln12a10 0.5
Kn3an12a11 Ln3a11 Ln12a11 0.5
Kn3an12a12 Ln3a12 Ln12a12 0.5
Kn3an12a13 Ln3a13 Ln12a13 0.5
Kn3an12a14 Ln3a14 Ln12a14 0.5
Kn3an12a15 Ln3a15 Ln12a15 0.5
Kn3an12a16 Ln3a16 Ln12a16 0.5
Kn3anva1 Ln3a1 Lnva1 0.5
Kn3anva2 Ln3a2 Lnva2 0.5
Kn3anva3 Ln3a3 Lnva3 0.5
Kn3anva4 Ln3a4 Lnva4 0.5
Kn3anva5 Ln3a5 Lnva5 0.5
Kn3anva6 Ln3a6 Lnva6 0.5
Kn3anva7 Ln3a7 Lnva7 0.5
Kn3anva8 Ln3a8 Lnva8 0.5
Kn3anva9 Ln3a9 Lnva9 0.5
Kn3anva10 Ln3a10 Lnva10 0.5
Kn3anva11 Ln3a11 Lnva11 0.5
Kn3anva12 Ln3a12 Lnva12 0.5
Kn3anva13 Ln3a13 Lnva13 0.5
Kn3anva14 Ln3a14 Lnva14 0.5
Kn3anva15 Ln3a15 Lnva15 0.5
Kn3anva16 Ln3a16 Lnva16 0.5
Kn4an5a1 Ln4a1 Ln5a1 0.8
Kn4an5a2 Ln4a2 Ln5a2 0.8
Kn4an5a3 Ln4a3 Ln5a3 0.8
Kn4an5a4 Ln4a4 Ln5a4 0.8
Kn4an5a5 Ln4a5 Ln5a5 0.8
Kn4an5a6 Ln4a6 Ln5a6 0.8
Kn4an5a7 Ln4a7 Ln5a7 0.8
Kn4an5a8 Ln4a8 Ln5a8 0.8
Kn4an5a9 Ln4a9 Ln5a9 0.8
Kn4an5a10 Ln4a10 Ln5a10 0.8
Kn4an5a11 Ln4a11 Ln5a11 0.8
Kn4an5a12 Ln4a12 Ln5a12 0.8
Kn4an5a13 Ln4a13 Ln5a13 0.8
Kn4an5a14 Ln4a14 Ln5a14 0.8
Kn4an5a15 Ln4a15 Ln5a15 0.8
Kn4an5a16 Ln4a16 Ln5a16 0.8
Kn4an6a1 Ln4a1 Ln6a1 0.7
Kn4an6a2 Ln4a2 Ln6a2 0.7
Kn4an6a3 Ln4a3 Ln6a3 0.7
Kn4an6a4 Ln4a4 Ln6a4 0.7
Kn4an6a5 Ln4a5 Ln6a5 0.7
Kn4an6a6 Ln4a6 Ln6a6 0.7
Kn4an6a7 Ln4a7 Ln6a7 0.7
Kn4an6a8 Ln4a8 Ln6a8 0.7
Kn4an6a9 Ln4a9 Ln6a9 0.7
Kn4an6a10 Ln4a10 Ln6a10 0.7
Kn4an6a11 Ln4a11 Ln6a11 0.7
Kn4an6a12 Ln4a12 Ln6a12 0.7
Kn4an6a13 Ln4a13 Ln6a13 0.7
Kn4an6a14 Ln4a14 Ln6a14 0.7
Kn4an6a15 Ln4a15 Ln6a15 0.7
Kn4an6a16 Ln4a16 Ln6a16 0.7
Kn4an7a1 Ln4a1 Ln7a1 0.7
Kn4an7a2 Ln4a2 Ln7a2 0.7
Kn4an7a3 Ln4a3 Ln7a3 0.7
Kn4an7a4 Ln4a4 Ln7a4 0.7
Kn4an7a5 Ln4a5 Ln7a5 0.7
Kn4an7a6 Ln4a6 Ln7a6 0.7
Kn4an7a7 Ln4a7 Ln7a7 0.7
Kn4an7a8 Ln4a8 Ln7a8 0.7
Kn4an7a9 Ln4a9 Ln7a9 0.7
Kn4an7a10 Ln4a10 Ln7a10 0.7
Kn4an7a11 Ln4a11 Ln7a11 0.7
Kn4an7a12 Ln4a12 Ln7a12 0.7
Kn4an7a13 Ln4a13 Ln7a13 0.7
Kn4an7a14 Ln4a14 Ln7a14 0.7
Kn4an7a15 Ln4a15 Ln7a15 0.7
Kn4an7a16 Ln4a16 Ln7a16 0.7
Kn4an8a1 Ln4a1 Ln8a1 0.6
Kn4an8a2 Ln4a2 Ln8a2 0.6
Kn4an8a3 Ln4a3 Ln8a3 0.6
Kn4an8a4 Ln4a4 Ln8a4 0.6
Kn4an8a5 Ln4a5 Ln8a5 0.6
Kn4an8a6 Ln4a6 Ln8a6 0.6
Kn4an8a7 Ln4a7 Ln8a7 0.6
Kn4an8a8 Ln4a8 Ln8a8 0.6
Kn4an8a9 Ln4a9 Ln8a9 0.6
Kn4an8a10 Ln4a10 Ln8a10 0.6
Kn4an8a11 Ln4a11 Ln8a11 0.6
Kn4an8a12 Ln4a12 Ln8a12 0.6
Kn4an8a13 Ln4a13 Ln8a13 0.6
Kn4an8a14 Ln4a14 Ln8a14 0.6
Kn4an8a15 Ln4a15 Ln8a15 0.6
Kn4an8a16 Ln4a16 Ln8a16 0.6
Kn4an9a1 Ln4a1 Ln9a1 0.6
Kn4an9a2 Ln4a2 Ln9a2 0.6
Kn4an9a3 Ln4a3 Ln9a3 0.6
Kn4an9a4 Ln4a4 Ln9a4 0.6
Kn4an9a5 Ln4a5 Ln9a5 0.6
Kn4an9a6 Ln4a6 Ln9a6 0.6
Kn4an9a7 Ln4a7 Ln9a7 0.6
Kn4an9a8 Ln4a8 Ln9a8 0.6
Kn4an9a9 Ln4a9 Ln9a9 0.6
Kn4an9a10 Ln4a10 Ln9a10 0.6
Kn4an9a11 Ln4a11 Ln9a11 0.6
Kn4an9a12 Ln4a12 Ln9a12 0.6
Kn4an9a13 Ln4a13 Ln9a13 0.6
Kn4an9a14 Ln4a14 Ln9a14 0.6
Kn4an9a15 Ln4a15 Ln9a15 0.6
Kn4an9a16 Ln4a16 Ln9a16 0.6
Kn4an10a1 Ln4a1 Ln10a1 0.6
Kn4an10a2 Ln4a2 Ln10a2 0.6
Kn4an10a3 Ln4a3 Ln10a3 0.6
Kn4an10a4 Ln4a4 Ln10a4 0.6
Kn4an10a5 Ln4a5 Ln10a5 0.6
Kn4an10a6 Ln4a6 Ln10a6 0.6
Kn4an10a7 Ln4a7 Ln10a7 0.6
Kn4an10a8 Ln4a8 Ln10a8 0.6
Kn4an10a9 Ln4a9 Ln10a9 0.6
Kn4an10a10 Ln4a10 Ln10a10 0.6
Kn4an10a11 Ln4a11 Ln10a11 0.6
Kn4an10a12 Ln4a12 Ln10a12 0.6
Kn4an10a13 Ln4a13 Ln10a13 0.6
Kn4an10a14 Ln4a14 Ln10a14 0.6
Kn4an10a15 Ln4a15 Ln10a15 0.6
Kn4an10a16 Ln4a16 Ln10a16 0.6
Kn4an11a1 Ln4a1 Ln11a1 0.6
Kn4an11a2 Ln4a2 Ln11a2 0.6
Kn4an11a3 Ln4a3 Ln11a3 0.6
Kn4an11a4 Ln4a4 Ln11a4 0.6
Kn4an11a5 Ln4a5 Ln11a5 0.6
Kn4an11a6 Ln4a6 Ln11a6 0.6
Kn4an11a7 Ln4a7 Ln11a7 0.6
Kn4an11a8 Ln4a8 Ln11a8 0.6
Kn4an11a9 Ln4a9 Ln11a9 0.6
Kn4an11a10 Ln4a10 Ln11a10 0.6
Kn4an11a11 Ln4a11 Ln11a11 0.6
Kn4an11a12 Ln4a12 Ln11a12 0.6
Kn4an11a13 Ln4a13 Ln11a13 0.6
Kn4an11a14 Ln4a14 Ln11a14 0.6
Kn4an11a15 Ln4a15 Ln11a15 0.6
Kn4an11a16 Ln4a16 Ln11a16 0.6
Kn4an12a1 Ln4a1 Ln12a1 0.6
Kn4an12a2 Ln4a2 Ln12a2 0.6
Kn4an12a3 Ln4a3 Ln12a3 0.6
Kn4an12a4 Ln4a4 Ln12a4 0.6
Kn4an12a5 Ln4a5 Ln12a5 0.6
Kn4an12a6 Ln4a6 Ln12a6 0.6
Kn4an12a7 Ln4a7 Ln12a7 0.6
Kn4an12a8 Ln4a8 Ln12a8 0.6
Kn4an12a9 Ln4a9 Ln12a9 0.6
Kn4an12a10 Ln4a10 Ln12a10 0.6
Kn4an12a11 Ln4a11 Ln12a11 0.6
Kn4an12a12 Ln4a12 Ln12a12 0.6
Kn4an12a13 Ln4a13 Ln12a13 0.6
Kn4an12a14 Ln4a14 Ln12a14 0.6
Kn4an12a15 Ln4a15 Ln12a15 0.6
Kn4an12a16 Ln4a16 Ln12a16 0.6
Kn4anva1 Ln4a1 Lnva1 0.5
Kn4anva2 Ln4a2 Lnva2 0.5
Kn4anva3 Ln4a3 Lnva3 0.5
Kn4anva4 Ln4a4 Lnva4 0.5
Kn4anva5 Ln4a5 Lnva5 0.5
Kn4anva6 Ln4a6 Lnva6 0.5
Kn4anva7 Ln4a7 Lnva7 0.5
Kn4anva8 Ln4a8 Lnva8 0.5
Kn4anva9 Ln4a9 Lnva9 0.5
Kn4anva10 Ln4a10 Lnva10 0.5
Kn4anva11 Ln4a11 Lnva11 0.5
Kn4anva12 Ln4a12 Lnva12 0.5
Kn4anva13 Ln4a13 Lnva13 0.5
Kn4anva14 Ln4a14 Lnva14 0.5
Kn4anva15 Ln4a15 Lnva15 0.5
Kn4anva16 Ln4a16 Lnva16 0.5
Kn5an6a1 Ln5a1 Ln6a1 0.8
Kn5an6a2 Ln5a2 Ln6a2 0.8
Kn5an6a3 Ln5a3 Ln6a3 0.8
Kn5an6a4 Ln5a4 Ln6a4 0.8
Kn5an6a5 Ln5a5 Ln6a5 0.8
Kn5an6a6 Ln5a6 Ln6a6 0.8
Kn5an6a7 Ln5a7 Ln6a7 0.8
Kn5an6a8 Ln5a8 Ln6a8 0.8
Kn5an6a9 Ln5a9 Ln6a9 0.8
Kn5an6a10 Ln5a10 Ln6a10 0.8
Kn5an6a11 Ln5a11 Ln6a11 0.8
Kn5an6a12 Ln5a12 Ln6a12 0.8
Kn5an6a13 Ln5a13 Ln6a13 0.8
Kn5an6a14 Ln5a14 Ln6a14 0.8
Kn5an6a15 Ln5a15 Ln6a15 0.8
Kn5an6a16 Ln5a16 Ln6a16 0.8
Kn5an7a1 Ln5a1 Ln7a1 0.7
Kn5an7a2 Ln5a2 Ln7a2 0.7
Kn5an7a3 Ln5a3 Ln7a3 0.7
Kn5an7a4 Ln5a4 Ln7a4 0.7
Kn5an7a5 Ln5a5 Ln7a5 0.7
Kn5an7a6 Ln5a6 Ln7a6 0.7
Kn5an7a7 Ln5a7 Ln7a7 0.7
Kn5an7a8 Ln5a8 Ln7a8 0.7
Kn5an7a9 Ln5a9 Ln7a9 0.7
Kn5an7a10 Ln5a10 Ln7a10 0.7
Kn5an7a11 Ln5a11 Ln7a11 0.7
Kn5an7a12 Ln5a12 Ln7a12 0.7
Kn5an7a13 Ln5a13 Ln7a13 0.7
Kn5an7a14 Ln5a14 Ln7a14 0.7
Kn5an7a15 Ln5a15 Ln7a15 0.7
Kn5an7a16 Ln5a16 Ln7a16 0.7
Kn5an8a1 Ln5a1 Ln8a1 0.7
Kn5an8a2 Ln5a2 Ln8a2 0.7
Kn5an8a3 Ln5a3 Ln8a3 0.7
Kn5an8a4 Ln5a4 Ln8a4 0.7
Kn5an8a5 Ln5a5 Ln8a5 0.7
Kn5an8a6 Ln5a6 Ln8a6 0.7
Kn5an8a7 Ln5a7 Ln8a7 0.7
Kn5an8a8 Ln5a8 Ln8a8 0.7
Kn5an8a9 Ln5a9 Ln8a9 0.7
Kn5an8a10 Ln5a10 Ln8a10 0.7
Kn5an8a11 Ln5a11 Ln8a11 0.7
Kn5an8a12 Ln5a12 Ln8a12 0.7
Kn5an8a13 Ln5a13 Ln8a13 0.7
Kn5an8a14 Ln5a14 Ln8a14 0.7
Kn5an8a15 Ln5a15 Ln8a15 0.7
Kn5an8a16 Ln5a16 Ln8a16 0.7
Kn5an9a1 Ln5a1 Ln9a1 0.6
Kn5an9a2 Ln5a2 Ln9a2 0.6
Kn5an9a3 Ln5a3 Ln9a3 0.6
Kn5an9a4 Ln5a4 Ln9a4 0.6
Kn5an9a5 Ln5a5 Ln9a5 0.6
Kn5an9a6 Ln5a6 Ln9a6 0.6
Kn5an9a7 Ln5a7 Ln9a7 0.6
Kn5an9a8 Ln5a8 Ln9a8 0.6
Kn5an9a9 Ln5a9 Ln9a9 0.6
Kn5an9a10 Ln5a10 Ln9a10 0.6
Kn5an9a11 Ln5a11 Ln9a11 0.6
Kn5an9a12 Ln5a12 Ln9a12 0.6
Kn5an9a13 Ln5a13 Ln9a13 0.6
Kn5an9a14 Ln5a14 Ln9a14 0.6
Kn5an9a15 Ln5a15 Ln9a15 0.6
Kn5an9a16 Ln5a16 Ln9a16 0.6
Kn5an10a1 Ln5a1 Ln10a1 0.6
Kn5an10a2 Ln5a2 Ln10a2 0.6
Kn5an10a3 Ln5a3 Ln10a3 0.6
Kn5an10a4 Ln5a4 Ln10a4 0.6
Kn5an10a5 Ln5a5 Ln10a5 0.6
Kn5an10a6 Ln5a6 Ln10a6 0.6
Kn5an10a7 Ln5a7 Ln10a7 0.6
Kn5an10a8 Ln5a8 Ln10a8 0.6
Kn5an10a9 Ln5a9 Ln10a9 0.6
Kn5an10a10 Ln5a10 Ln10a10 0.6
Kn5an10a11 Ln5a11 Ln10a11 0.6
Kn5an10a12 Ln5a12 Ln10a12 0.6
Kn5an10a13 Ln5a13 Ln10a13 0.6
Kn5an10a14 Ln5a14 Ln10a14 0.6
Kn5an10a15 Ln5a15 Ln10a15 0.6
Kn5an10a16 Ln5a16 Ln10a16 0.6
Kn5an11a1 Ln5a1 Ln11a1 0.6
Kn5an11a2 Ln5a2 Ln11a2 0.6
Kn5an11a3 Ln5a3 Ln11a3 0.6
Kn5an11a4 Ln5a4 Ln11a4 0.6
Kn5an11a5 Ln5a5 Ln11a5 0.6
Kn5an11a6 Ln5a6 Ln11a6 0.6
Kn5an11a7 Ln5a7 Ln11a7 0.6
Kn5an11a8 Ln5a8 Ln11a8 0.6
Kn5an11a9 Ln5a9 Ln11a9 0.6
Kn5an11a10 Ln5a10 Ln11a10 0.6
Kn5an11a11 Ln5a11 Ln11a11 0.6
Kn5an11a12 Ln5a12 Ln11a12 0.6
Kn5an11a13 Ln5a13 Ln11a13 0.6
Kn5an11a14 Ln5a14 Ln11a14 0.6
Kn5an11a15 Ln5a15 Ln11a15 0.6
Kn5an11a16 Ln5a16 Ln11a16 0.6
Kn5an12a1 Ln5a1 Ln12a1 0.6
Kn5an12a2 Ln5a2 Ln12a2 0.6
Kn5an12a3 Ln5a3 Ln12a3 0.6
Kn5an12a4 Ln5a4 Ln12a4 0.6
Kn5an12a5 Ln5a5 Ln12a5 0.6
Kn5an12a6 Ln5a6 Ln12a6 0.6
Kn5an12a7 Ln5a7 Ln12a7 0.6
Kn5an12a8 Ln5a8 Ln12a8 0.6
Kn5an12a9 Ln5a9 Ln12a9 0.6
Kn5an12a10 Ln5a10 Ln12a10 0.6
Kn5an12a11 Ln5a11 Ln12a11 0.6
Kn5an12a12 Ln5a12 Ln12a12 0.6
Kn5an12a13 Ln5a13 Ln12a13 0.6
Kn5an12a14 Ln5a14 Ln12a14 0.6
Kn5an12a15 Ln5a15 Ln12a15 0.6
Kn5an12a16 Ln5a16 Ln12a16 0.6
Kn5anva1 Ln5a1 Lnva1 0.6
Kn5anva2 Ln5a2 Lnva2 0.6
Kn5anva3 Ln5a3 Lnva3 0.6
Kn5anva4 Ln5a4 Lnva4 0.6
Kn5anva5 Ln5a5 Lnva5 0.6
Kn5anva6 Ln5a6 Lnva6 0.6
Kn5anva7 Ln5a7 Lnva7 0.6
Kn5anva8 Ln5a8 Lnva8 0.6
Kn5anva9 Ln5a9 Lnva9 0.6
Kn5anva10 Ln5a10 Lnva10 0.6
Kn5anva11 Ln5a11 Lnva11 0.6
Kn5anva12 Ln5a12 Lnva12 0.6
Kn5anva13 Ln5a13 Lnva13 0.6
Kn5anva14 Ln5a14 Lnva14 0.6
Kn5anva15 Ln5a15 Lnva15 0.6
Kn5anva16 Ln5a16 Lnva16 0.6
Kn6an7a1 Ln6a1 Ln7a1 0.8
Kn6an7a2 Ln6a2 Ln7a2 0.8
Kn6an7a3 Ln6a3 Ln7a3 0.8
Kn6an7a4 Ln6a4 Ln7a4 0.8
Kn6an7a5 Ln6a5 Ln7a5 0.8
Kn6an7a6 Ln6a6 Ln7a6 0.8
Kn6an7a7 Ln6a7 Ln7a7 0.8
Kn6an7a8 Ln6a8 Ln7a8 0.8
Kn6an7a9 Ln6a9 Ln7a9 0.8
Kn6an7a10 Ln6a10 Ln7a10 0.8
Kn6an7a11 Ln6a11 Ln7a11 0.8
Kn6an7a12 Ln6a12 Ln7a12 0.8
Kn6an7a13 Ln6a13 Ln7a13 0.8
Kn6an7a14 Ln6a14 Ln7a14 0.8
Kn6an7a15 Ln6a15 Ln7a15 0.8
Kn6an7a16 Ln6a16 Ln7a16 0.8
Kn6an8a1 Ln6a1 Ln8a1 0.7
Kn6an8a2 Ln6a2 Ln8a2 0.7
Kn6an8a3 Ln6a3 Ln8a3 0.7
Kn6an8a4 Ln6a4 Ln8a4 0.7
Kn6an8a5 Ln6a5 Ln8a5 0.7
Kn6an8a6 Ln6a6 Ln8a6 0.7
Kn6an8a7 Ln6a7 Ln8a7 0.7
Kn6an8a8 Ln6a8 Ln8a8 0.7
Kn6an8a9 Ln6a9 Ln8a9 0.7
Kn6an8a10 Ln6a10 Ln8a10 0.7
Kn6an8a11 Ln6a11 Ln8a11 0.7
Kn6an8a12 Ln6a12 Ln8a12 0.7
Kn6an8a13 Ln6a13 Ln8a13 0.7
Kn6an8a14 Ln6a14 Ln8a14 0.7
Kn6an8a15 Ln6a15 Ln8a15 0.7
Kn6an8a16 Ln6a16 Ln8a16 0.7
Kn6an9a1 Ln6a1 Ln9a1 0.7
Kn6an9a2 Ln6a2 Ln9a2 0.7
Kn6an9a3 Ln6a3 Ln9a3 0.7
Kn6an9a4 Ln6a4 Ln9a4 0.7
Kn6an9a5 Ln6a5 Ln9a5 0.7
Kn6an9a6 Ln6a6 Ln9a6 0.7
Kn6an9a7 Ln6a7 Ln9a7 0.7
Kn6an9a8 Ln6a8 Ln9a8 0.7
Kn6an9a9 Ln6a9 Ln9a9 0.7
Kn6an9a10 Ln6a10 Ln9a10 0.7
Kn6an9a11 Ln6a11 Ln9a11 0.7
Kn6an9a12 Ln6a12 Ln9a12 0.7
Kn6an9a13 Ln6a13 Ln9a13 0.7
Kn6an9a14 Ln6a14 Ln9a14 0.7
Kn6an9a15 Ln6a15 Ln9a15 0.7
Kn6an9a16 Ln6a16 Ln9a16 0.7
Kn6an10a1 Ln6a1 Ln10a1 0.6
Kn6an10a2 Ln6a2 Ln10a2 0.6
Kn6an10a3 Ln6a3 Ln10a3 0.6
Kn6an10a4 Ln6a4 Ln10a4 0.6
Kn6an10a5 Ln6a5 Ln10a5 0.6
Kn6an10a6 Ln6a6 Ln10a6 0.6
Kn6an10a7 Ln6a7 Ln10a7 0.6
Kn6an10a8 Ln6a8 Ln10a8 0.6
Kn6an10a9 Ln6a9 Ln10a9 0.6
Kn6an10a10 Ln6a10 Ln10a10 0.6
Kn6an10a11 Ln6a11 Ln10a11 0.6
Kn6an10a12 Ln6a12 Ln10a12 0.6
Kn6an10a13 Ln6a13 Ln10a13 0.6
Kn6an10a14 Ln6a14 Ln10a14 0.6
Kn6an10a15 Ln6a15 Ln10a15 0.6
Kn6an10a16 Ln6a16 Ln10a16 0.6
Kn6an11a1 Ln6a1 Ln11a1 0.6
Kn6an11a2 Ln6a2 Ln11a2 0.6
Kn6an11a3 Ln6a3 Ln11a3 0.6
Kn6an11a4 Ln6a4 Ln11a4 0.6
Kn6an11a5 Ln6a5 Ln11a5 0.6
Kn6an11a6 Ln6a6 Ln11a6 0.6
Kn6an11a7 Ln6a7 Ln11a7 0.6
Kn6an11a8 Ln6a8 Ln11a8 0.6
Kn6an11a9 Ln6a9 Ln11a9 0.6
Kn6an11a10 Ln6a10 Ln11a10 0.6
Kn6an11a11 Ln6a11 Ln11a11 0.6
Kn6an11a12 Ln6a12 Ln11a12 0.6
Kn6an11a13 Ln6a13 Ln11a13 0.6
Kn6an11a14 Ln6a14 Ln11a14 0.6
Kn6an11a15 Ln6a15 Ln11a15 0.6
Kn6an11a16 Ln6a16 Ln11a16 0.6
Kn6an12a1 Ln6a1 Ln12a1 0.6
Kn6an12a2 Ln6a2 Ln12a2 0.6
Kn6an12a3 Ln6a3 Ln12a3 0.6
Kn6an12a4 Ln6a4 Ln12a4 0.6
Kn6an12a5 Ln6a5 Ln12a5 0.6
Kn6an12a6 Ln6a6 Ln12a6 0.6
Kn6an12a7 Ln6a7 Ln12a7 0.6
Kn6an12a8 Ln6a8 Ln12a8 0.6
Kn6an12a9 Ln6a9 Ln12a9 0.6
Kn6an12a10 Ln6a10 Ln12a10 0.6
Kn6an12a11 Ln6a11 Ln12a11 0.6
Kn6an12a12 Ln6a12 Ln12a12 0.6
Kn6an12a13 Ln6a13 Ln12a13 0.6
Kn6an12a14 Ln6a14 Ln12a14 0.6
Kn6an12a15 Ln6a15 Ln12a15 0.6
Kn6an12a16 Ln6a16 Ln12a16 0.6
Kn6anva1 Ln6a1 Lnva1 0.6
Kn6anva2 Ln6a2 Lnva2 0.6
Kn6anva3 Ln6a3 Lnva3 0.6
Kn6anva4 Ln6a4 Lnva4 0.6
Kn6anva5 Ln6a5 Lnva5 0.6
Kn6anva6 Ln6a6 Lnva6 0.6
Kn6anva7 Ln6a7 Lnva7 0.6
Kn6anva8 Ln6a8 Lnva8 0.6
Kn6anva9 Ln6a9 Lnva9 0.6
Kn6anva10 Ln6a10 Lnva10 0.6
Kn6anva11 Ln6a11 Lnva11 0.6
Kn6anva12 Ln6a12 Lnva12 0.6
Kn6anva13 Ln6a13 Lnva13 0.6
Kn6anva14 Ln6a14 Lnva14 0.6
Kn6anva15 Ln6a15 Lnva15 0.6
Kn6anva16 Ln6a16 Lnva16 0.6
Kn7an8a1 Ln7a1 Ln8a1 0.8
Kn7an8a2 Ln7a2 Ln8a2 0.8
Kn7an8a3 Ln7a3 Ln8a3 0.8
Kn7an8a4 Ln7a4 Ln8a4 0.8
Kn7an8a5 Ln7a5 Ln8a5 0.8
Kn7an8a6 Ln7a6 Ln8a6 0.8
Kn7an8a7 Ln7a7 Ln8a7 0.8
Kn7an8a8 Ln7a8 Ln8a8 0.8
Kn7an8a9 Ln7a9 Ln8a9 0.8
Kn7an8a10 Ln7a10 Ln8a10 0.8
Kn7an8a11 Ln7a11 Ln8a11 0.8
Kn7an8a12 Ln7a12 Ln8a12 0.8
Kn7an8a13 Ln7a13 Ln8a13 0.8
Kn7an8a14 Ln7a14 Ln8a14 0.8
Kn7an8a15 Ln7a15 Ln8a15 0.8
Kn7an8a16 Ln7a16 Ln8a16 0.8
Kn7an9a1 Ln7a1 Ln9a1 0.7
Kn7an9a2 Ln7a2 Ln9a2 0.7
Kn7an9a3 Ln7a3 Ln9a3 0.7
Kn7an9a4 Ln7a4 Ln9a4 0.7
Kn7an9a5 Ln7a5 Ln9a5 0.7
Kn7an9a6 Ln7a6 Ln9a6 0.7
Kn7an9a7 Ln7a7 Ln9a7 0.7
Kn7an9a8 Ln7a8 Ln9a8 0.7
Kn7an9a9 Ln7a9 Ln9a9 0.7
Kn7an9a10 Ln7a10 Ln9a10 0.7
Kn7an9a11 Ln7a11 Ln9a11 0.7
Kn7an9a12 Ln7a12 Ln9a12 0.7
Kn7an9a13 Ln7a13 Ln9a13 0.7
Kn7an9a14 Ln7a14 Ln9a14 0.7
Kn7an9a15 Ln7a15 Ln9a15 0.7
Kn7an9a16 Ln7a16 Ln9a16 0.7
Kn7an10a1 Ln7a1 Ln10a1 0.7
Kn7an10a2 Ln7a2 Ln10a2 0.7
Kn7an10a3 Ln7a3 Ln10a3 0.7
Kn7an10a4 Ln7a4 Ln10a4 0.7
Kn7an10a5 Ln7a5 Ln10a5 0.7
Kn7an10a6 Ln7a6 Ln10a6 0.7
Kn7an10a7 Ln7a7 Ln10a7 0.7
Kn7an10a8 Ln7a8 Ln10a8 0.7
Kn7an10a9 Ln7a9 Ln10a9 0.7
Kn7an10a10 Ln7a10 Ln10a10 0.7
Kn7an10a11 Ln7a11 Ln10a11 0.7
Kn7an10a12 Ln7a12 Ln10a12 0.7
Kn7an10a13 Ln7a13 Ln10a13 0.7
Kn7an10a14 Ln7a14 Ln10a14 0.7
Kn7an10a15 Ln7a15 Ln10a15 0.7
Kn7an10a16 Ln7a16 Ln10a16 0.7
Kn7an11a1 Ln7a1 Ln11a1 0.6
Kn7an11a2 Ln7a2 Ln11a2 0.6
Kn7an11a3 Ln7a3 Ln11a3 0.6
Kn7an11a4 Ln7a4 Ln11a4 0.6
Kn7an11a5 Ln7a5 Ln11a5 0.6
Kn7an11a6 Ln7a6 Ln11a6 0.6
Kn7an11a7 Ln7a7 Ln11a7 0.6
Kn7an11a8 Ln7a8 Ln11a8 0.6
Kn7an11a9 Ln7a9 Ln11a9 0.6
Kn7an11a10 Ln7a10 Ln11a10 0.6
Kn7an11a11 Ln7a11 Ln11a11 0.6
Kn7an11a12 Ln7a12 Ln11a12 0.6
Kn7an11a13 Ln7a13 Ln11a13 0.6
Kn7an11a14 Ln7a14 Ln11a14 0.6
Kn7an11a15 Ln7a15 Ln11a15 0.6
Kn7an11a16 Ln7a16 Ln11a16 0.6
Kn7an12a1 Ln7a1 Ln12a1 0.6
Kn7an12a2 Ln7a2 Ln12a2 0.6
Kn7an12a3 Ln7a3 Ln12a3 0.6
Kn7an12a4 Ln7a4 Ln12a4 0.6
Kn7an12a5 Ln7a5 Ln12a5 0.6
Kn7an12a6 Ln7a6 Ln12a6 0.6
Kn7an12a7 Ln7a7 Ln12a7 0.6
Kn7an12a8 Ln7a8 Ln12a8 0.6
Kn7an12a9 Ln7a9 Ln12a9 0.6
Kn7an12a10 Ln7a10 Ln12a10 0.6
Kn7an12a11 Ln7a11 Ln12a11 0.6
Kn7an12a12 Ln7a12 Ln12a12 0.6
Kn7an12a13 Ln7a13 Ln12a13 0.6
Kn7an12a14 Ln7a14 Ln12a14 0.6
Kn7an12a15 Ln7a15 Ln12a15 0.6
Kn7an12a16 Ln7a16 Ln12a16 0.6
Kn7anva1 Ln7a1 Lnva1 0.6
Kn7anva2 Ln7a2 Lnva2 0.6
Kn7anva3 Ln7a3 Lnva3 0.6
Kn7anva4 Ln7a4 Lnva4 0.6
Kn7anva5 Ln7a5 Lnva5 0.6
Kn7anva6 Ln7a6 Lnva6 0.6
Kn7anva7 Ln7a7 Lnva7 0.6
Kn7anva8 Ln7a8 Lnva8 0.6
Kn7anva9 Ln7a9 Lnva9 0.6
Kn7anva10 Ln7a10 Lnva10 0.6
Kn7anva11 Ln7a11 Lnva11 0.6
Kn7anva12 Ln7a12 Lnva12 0.6
Kn7anva13 Ln7a13 Lnva13 0.6
Kn7anva14 Ln7a14 Lnva14 0.6
Kn7anva15 Ln7a15 Lnva15 0.6
Kn7anva16 Ln7a16 Lnva16 0.6
Kn8an9a1 Ln8a1 Ln9a1 0.8
Kn8an9a2 Ln8a2 Ln9a2 0.8
Kn8an9a3 Ln8a3 Ln9a3 0.8
Kn8an9a4 Ln8a4 Ln9a4 0.8
Kn8an9a5 Ln8a5 Ln9a5 0.8
Kn8an9a6 Ln8a6 Ln9a6 0.8
Kn8an9a7 Ln8a7 Ln9a7 0.8
Kn8an9a8 Ln8a8 Ln9a8 0.8
Kn8an9a9 Ln8a9 Ln9a9 0.8
Kn8an9a10 Ln8a10 Ln9a10 0.8
Kn8an9a11 Ln8a11 Ln9a11 0.8
Kn8an9a12 Ln8a12 Ln9a12 0.8
Kn8an9a13 Ln8a13 Ln9a13 0.8
Kn8an9a14 Ln8a14 Ln9a14 0.8
Kn8an9a15 Ln8a15 Ln9a15 0.8
Kn8an9a16 Ln8a16 Ln9a16 0.8
Kn8an10a1 Ln8a1 Ln10a1 0.7
Kn8an10a2 Ln8a2 Ln10a2 0.7
Kn8an10a3 Ln8a3 Ln10a3 0.7
Kn8an10a4 Ln8a4 Ln10a4 0.7
Kn8an10a5 Ln8a5 Ln10a5 0.7
Kn8an10a6 Ln8a6 Ln10a6 0.7
Kn8an10a7 Ln8a7 Ln10a7 0.7
Kn8an10a8 Ln8a8 Ln10a8 0.7
Kn8an10a9 Ln8a9 Ln10a9 0.7
Kn8an10a10 Ln8a10 Ln10a10 0.7
Kn8an10a11 Ln8a11 Ln10a11 0.7
Kn8an10a12 Ln8a12 Ln10a12 0.7
Kn8an10a13 Ln8a13 Ln10a13 0.7
Kn8an10a14 Ln8a14 Ln10a14 0.7
Kn8an10a15 Ln8a15 Ln10a15 0.7
Kn8an10a16 Ln8a16 Ln10a16 0.7
Kn8an11a1 Ln8a1 Ln11a1 0.7
Kn8an11a2 Ln8a2 Ln11a2 0.7
Kn8an11a3 Ln8a3 Ln11a3 0.7
Kn8an11a4 Ln8a4 Ln11a4 0.7
Kn8an11a5 Ln8a5 Ln11a5 0.7
Kn8an11a6 Ln8a6 Ln11a6 0.7
Kn8an11a7 Ln8a7 Ln11a7 0.7
Kn8an11a8 Ln8a8 Ln11a8 0.7
Kn8an11a9 Ln8a9 Ln11a9 0.7
Kn8an11a10 Ln8a10 Ln11a10 0.7
Kn8an11a11 Ln8a11 Ln11a11 0.7
Kn8an11a12 Ln8a12 Ln11a12 0.7
Kn8an11a13 Ln8a13 Ln11a13 0.7
Kn8an11a14 Ln8a14 Ln11a14 0.7
Kn8an11a15 Ln8a15 Ln11a15 0.7
Kn8an11a16 Ln8a16 Ln11a16 0.7
Kn8an12a1 Ln8a1 Ln12a1 0.6
Kn8an12a2 Ln8a2 Ln12a2 0.6
Kn8an12a3 Ln8a3 Ln12a3 0.6
Kn8an12a4 Ln8a4 Ln12a4 0.6
Kn8an12a5 Ln8a5 Ln12a5 0.6
Kn8an12a6 Ln8a6 Ln12a6 0.6
Kn8an12a7 Ln8a7 Ln12a7 0.6
Kn8an12a8 Ln8a8 Ln12a8 0.6
Kn8an12a9 Ln8a9 Ln12a9 0.6
Kn8an12a10 Ln8a10 Ln12a10 0.6
Kn8an12a11 Ln8a11 Ln12a11 0.6
Kn8an12a12 Ln8a12 Ln12a12 0.6
Kn8an12a13 Ln8a13 Ln12a13 0.6
Kn8an12a14 Ln8a14 Ln12a14 0.6
Kn8an12a15 Ln8a15 Ln12a15 0.6
Kn8an12a16 Ln8a16 Ln12a16 0.6
Kn8anva1 Ln8a1 Lnva1 0.6
Kn8anva2 Ln8a2 Lnva2 0.6
Kn8anva3 Ln8a3 Lnva3 0.6
Kn8anva4 Ln8a4 Lnva4 0.6
Kn8anva5 Ln8a5 Lnva5 0.6
Kn8anva6 Ln8a6 Lnva6 0.6
Kn8anva7 Ln8a7 Lnva7 0.6
Kn8anva8 Ln8a8 Lnva8 0.6
Kn8anva9 Ln8a9 Lnva9 0.6
Kn8anva10 Ln8a10 Lnva10 0.6
Kn8anva11 Ln8a11 Lnva11 0.6
Kn8anva12 Ln8a12 Lnva12 0.6
Kn8anva13 Ln8a13 Lnva13 0.6
Kn8anva14 Ln8a14 Lnva14 0.6
Kn8anva15 Ln8a15 Lnva15 0.6
Kn8anva16 Ln8a16 Lnva16 0.6
Kn9an10a1 Ln9a1 Ln10a1 0.8
Kn9an10a2 Ln9a2 Ln10a2 0.8
Kn9an10a3 Ln9a3 Ln10a3 0.8
Kn9an10a4 Ln9a4 Ln10a4 0.8
Kn9an10a5 Ln9a5 Ln10a5 0.8
Kn9an10a6 Ln9a6 Ln10a6 0.8
Kn9an10a7 Ln9a7 Ln10a7 0.8
Kn9an10a8 Ln9a8 Ln10a8 0.8
Kn9an10a9 Ln9a9 Ln10a9 0.8
Kn9an10a10 Ln9a10 Ln10a10 0.8
Kn9an10a11 Ln9a11 Ln10a11 0.8
Kn9an10a12 Ln9a12 Ln10a12 0.8
Kn9an10a13 Ln9a13 Ln10a13 0.8
Kn9an10a14 Ln9a14 Ln10a14 0.8
Kn9an10a15 Ln9a15 Ln10a15 0.8
Kn9an10a16 Ln9a16 Ln10a16 0.8
Kn9an11a1 Ln9a1 Ln11a1 0.7
Kn9an11a2 Ln9a2 Ln11a2 0.7
Kn9an11a3 Ln9a3 Ln11a3 0.7
Kn9an11a4 Ln9a4 Ln11a4 0.7
Kn9an11a5 Ln9a5 Ln11a5 0.7
Kn9an11a6 Ln9a6 Ln11a6 0.7
Kn9an11a7 Ln9a7 Ln11a7 0.7
Kn9an11a8 Ln9a8 Ln11a8 0.7
Kn9an11a9 Ln9a9 Ln11a9 0.7
Kn9an11a10 Ln9a10 Ln11a10 0.7
Kn9an11a11 Ln9a11 Ln11a11 0.7
Kn9an11a12 Ln9a12 Ln11a12 0.7
Kn9an11a13 Ln9a13 Ln11a13 0.7
Kn9an11a14 Ln9a14 Ln11a14 0.7
Kn9an11a15 Ln9a15 Ln11a15 0.7
Kn9an11a16 Ln9a16 Ln11a16 0.7
Kn9an12a1 Ln9a1 Ln12a1 0.7
Kn9an12a2 Ln9a2 Ln12a2 0.7
Kn9an12a3 Ln9a3 Ln12a3 0.7
Kn9an12a4 Ln9a4 Ln12a4 0.7
Kn9an12a5 Ln9a5 Ln12a5 0.7
Kn9an12a6 Ln9a6 Ln12a6 0.7
Kn9an12a7 Ln9a7 Ln12a7 0.7
Kn9an12a8 Ln9a8 Ln12a8 0.7
Kn9an12a9 Ln9a9 Ln12a9 0.7
Kn9an12a10 Ln9a10 Ln12a10 0.7
Kn9an12a11 Ln9a11 Ln12a11 0.7
Kn9an12a12 Ln9a12 Ln12a12 0.7
Kn9an12a13 Ln9a13 Ln12a13 0.7
Kn9an12a14 Ln9a14 Ln12a14 0.7
Kn9an12a15 Ln9a15 Ln12a15 0.7
Kn9an12a16 Ln9a16 Ln12a16 0.7
Kn9anva1 Ln9a1 Lnva1 0.6
Kn9anva2 Ln9a2 Lnva2 0.6
Kn9anva3 Ln9a3 Lnva3 0.6
Kn9anva4 Ln9a4 Lnva4 0.6
Kn9anva5 Ln9a5 Lnva5 0.6
Kn9anva6 Ln9a6 Lnva6 0.6
Kn9anva7 Ln9a7 Lnva7 0.6
Kn9anva8 Ln9a8 Lnva8 0.6
Kn9anva9 Ln9a9 Lnva9 0.6
Kn9anva10 Ln9a10 Lnva10 0.6
Kn9anva11 Ln9a11 Lnva11 0.6
Kn9anva12 Ln9a12 Lnva12 0.6
Kn9anva13 Ln9a13 Lnva13 0.6
Kn9anva14 Ln9a14 Lnva14 0.6
Kn9anva15 Ln9a15 Lnva15 0.6
Kn9anva16 Ln9a16 Lnva16 0.6
Kn10an11a1 Ln10a1 Ln11a1 0.8
Kn10an11a2 Ln10a2 Ln11a2 0.8
Kn10an11a3 Ln10a3 Ln11a3 0.8
Kn10an11a4 Ln10a4 Ln11a4 0.8
Kn10an11a5 Ln10a5 Ln11a5 0.8
Kn10an11a6 Ln10a6 Ln11a6 0.8
Kn10an11a7 Ln10a7 Ln11a7 0.8
Kn10an11a8 Ln10a8 Ln11a8 0.8
Kn10an11a9 Ln10a9 Ln11a9 0.8
Kn10an11a10 Ln10a10 Ln11a10 0.8
Kn10an11a11 Ln10a11 Ln11a11 0.8
Kn10an11a12 Ln10a12 Ln11a12 0.8
Kn10an11a13 Ln10a13 Ln11a13 0.8
Kn10an11a14 Ln10a14 Ln11a14 0.8
Kn10an11a15 Ln10a15 Ln11a15 0.8
Kn10an11a16 Ln10a16 Ln11a16 0.8
Kn10an12a1 Ln10a1 Ln12a1 0.7
Kn10an12a2 Ln10a2 Ln12a2 0.7
Kn10an12a3 Ln10a3 Ln12a3 0.7
Kn10an12a4 Ln10a4 Ln12a4 0.7
Kn10an12a5 Ln10a5 Ln12a5 0.7
Kn10an12a6 Ln10a6 Ln12a6 0.7
Kn10an12a7 Ln10a7 Ln12a7 0.7
Kn10an12a8 Ln10a8 Ln12a8 0.7
Kn10an12a9 Ln10a9 Ln12a9 0.7
Kn10an12a10 Ln10a10 Ln12a10 0.7
Kn10an12a11 Ln10a11 Ln12a11 0.7
Kn10an12a12 Ln10a12 Ln12a12 0.7
Kn10an12a13 Ln10a13 Ln12a13 0.7
Kn10an12a14 Ln10a14 Ln12a14 0.7
Kn10an12a15 Ln10a15 Ln12a15 0.7
Kn10an12a16 Ln10a16 Ln12a16 0.7
Kn10anva1 Ln10a1 Lnva1 0.7
Kn10anva2 Ln10a2 Lnva2 0.7
Kn10anva3 Ln10a3 Lnva3 0.7
Kn10anva4 Ln10a4 Lnva4 0.7
Kn10anva5 Ln10a5 Lnva5 0.7
Kn10anva6 Ln10a6 Lnva6 0.7
Kn10anva7 Ln10a7 Lnva7 0.7
Kn10anva8 Ln10a8 Lnva8 0.7
Kn10anva9 Ln10a9 Lnva9 0.7
Kn10anva10 Ln10a10 Lnva10 0.7
Kn10anva11 Ln10a11 Lnva11 0.7
Kn10anva12 Ln10a12 Lnva12 0.7
Kn10anva13 Ln10a13 Lnva13 0.7
Kn10anva14 Ln10a14 Lnva14 0.7
Kn10anva15 Ln10a15 Lnva15 0.7
Kn10anva16 Ln10a16 Lnva16 0.7
Kn11an12a1 Ln11a1 Ln12a1 0.8
Kn11an12a2 Ln11a2 Ln12a2 0.8
Kn11an12a3 Ln11a3 Ln12a3 0.8
Kn11an12a4 Ln11a4 Ln12a4 0.8
Kn11an12a5 Ln11a5 Ln12a5 0.8
Kn11an12a6 Ln11a6 Ln12a6 0.8
Kn11an12a7 Ln11a7 Ln12a7 0.8
Kn11an12a8 Ln11a8 Ln12a8 0.8
Kn11an12a9 Ln11a9 Ln12a9 0.8
Kn11an12a10 Ln11a10 Ln12a10 0.8
Kn11an12a11 Ln11a11 Ln12a11 0.8
Kn11an12a12 Ln11a12 Ln12a12 0.8
Kn11an12a13 Ln11a13 Ln12a13 0.8
Kn11an12a14 Ln11a14 Ln12a14 0.8
Kn11an12a15 Ln11a15 Ln12a15 0.8
Kn11an12a16 Ln11a16 Ln12a16 0.8
Kn11anva1 Ln11a1 Lnva1 0.7
Kn11anva2 Ln11a2 Lnva2 0.7
Kn11anva3 Ln11a3 Lnva3 0.7
Kn11anva4 Ln11a4 Lnva4 0.7
Kn11anva5 Ln11a5 Lnva5 0.7
Kn11anva6 Ln11a6 Lnva6 0.7
Kn11anva7 Ln11a7 Lnva7 0.7
Kn11anva8 Ln11a8 Lnva8 0.7
Kn11anva9 Ln11a9 Lnva9 0.7
Kn11anva10 Ln11a10 Lnva10 0.7
Kn11anva11 Ln11a11 Lnva11 0.7
Kn11anva12 Ln11a12 Lnva12 0.7
Kn11anva13 Ln11a13 Lnva13 0.7
Kn11anva14 Ln11a14 Lnva14 0.7
Kn11anva15 Ln11a15 Lnva15 0.7
Kn11anva16 Ln11a16 Lnva16 0.7
Kn12anva1 Ln12a1 Lnva1 0.8
Kn12anva2 Ln12a2 Lnva2 0.8
Kn12anva3 Ln12a3 Lnva3 0.8
Kn12anva4 Ln12a4 Lnva4 0.8
Kn12anva5 Ln12a5 Lnva5 0.8
Kn12anva6 Ln12a6 Lnva6 0.8
Kn12anva7 Ln12a7 Lnva7 0.8
Kn12anva8 Ln12a8 Lnva8 0.8
Kn12anva9 Ln12a9 Lnva9 0.8
Kn12anva10 Ln12a10 Lnva10 0.8
Kn12anva11 Ln12a11 Lnva11 0.8
Kn12anva12 Ln12a12 Lnva12 0.8
Kn12anva13 Ln12a13 Lnva13 0.8
Kn12anva14 Ln12a14 Lnva14 0.8
Kn12anva15 Ln12a15 Lnva15 0.8
Kn12anva16 Ln12a16 Lnva16 0.8
Cngan1a1 TDnga1 TDn1a1 2e-014
Cngan1a2 TDnga3 TDn1a3 3e-014
Cngan1a3 TDnga5 TDn1a5 3e-014
Cngan1a4 TDnga7 TDn1a7 3e-014
Cngan1a5 TDnga9 TDn1a9 3e-014
Cngan1a6 TDnga11 TDn1a11 3e-014
Cngan1a7 TDnga13 TDn1a13 3e-014
Cngan1a8 TDnga15 TDn1a15 3e-014
Cngan1a9 TDnga17 TDn1a17 3e-014
Cngan1a10 TDnga19 TDn1a19 3e-014
Cngan1a11 TDnga21 TDn1a21 3e-014
Cngan1a12 TDnga23 TDn1a23 3e-014
Cngan1a13 TDnga25 TDn1a25 3e-014
Cngan1a14 TDnga27 TDn1a27 3e-014
Cngan1a15 TDnga29 TDn1a29 3e-014
Cngan1a16 TDnga31 TDn1a31 3e-014
Cngan1a17 TDnga33 TDn1a33 2e-014
Cngan2a1 TDnga1 TDn2a1 7e-015
Cngan2a2 TDnga3 TDn2a3 1e-014
Cngan2a3 TDnga5 TDn2a5 1e-014
Cngan2a4 TDnga7 TDn2a7 1e-014
Cngan2a5 TDnga9 TDn2a9 1e-014
Cngan2a6 TDnga11 TDn2a11 1e-014
Cngan2a7 TDnga13 TDn2a13 1e-014
Cngan2a8 TDnga15 TDn2a15 1e-014
Cngan2a9 TDnga17 TDn2a17 1e-014
Cngan2a10 TDnga19 TDn2a19 1e-014
Cngan2a11 TDnga21 TDn2a21 1e-014
Cngan2a12 TDnga23 TDn2a23 1e-014
Cngan2a13 TDnga25 TDn2a25 1e-014
Cngan2a14 TDnga27 TDn2a27 1e-014
Cngan2a15 TDnga29 TDn2a29 1e-014
Cngan2a16 TDnga31 TDn2a31 1e-014
Cngan2a17 TDnga33 TDn2a33 7e-015
Cngan3a1 TDnga1 TDn3a1 6e-015
Cngan3a2 TDnga3 TDn3a3 1e-014
Cngan3a3 TDnga5 TDn3a5 1e-014
Cngan3a4 TDnga7 TDn3a7 1e-014
Cngan3a5 TDnga9 TDn3a9 1e-014
Cngan3a6 TDnga11 TDn3a11 1e-014
Cngan3a7 TDnga13 TDn3a13 1e-014
Cngan3a8 TDnga15 TDn3a15 1e-014
Cngan3a9 TDnga17 TDn3a17 1e-014
Cngan3a10 TDnga19 TDn3a19 1e-014
Cngan3a11 TDnga21 TDn3a21 1e-014
Cngan3a12 TDnga23 TDn3a23 1e-014
Cngan3a13 TDnga25 TDn3a25 1e-014
Cngan3a14 TDnga27 TDn3a27 1e-014
Cngan3a15 TDnga29 TDn3a29 1e-014
Cngan3a16 TDnga31 TDn3a31 1e-014
Cngan3a17 TDnga33 TDn3a33 6e-015
Cngan4a1 TDnga1 TDn4a1 6e-015
Cngan4a2 TDnga3 TDn4a3 1e-014
Cngan4a3 TDnga5 TDn4a5 1e-014
Cngan4a4 TDnga7 TDn4a7 1e-014
Cngan4a5 TDnga9 TDn4a9 1e-014
Cngan4a6 TDnga11 TDn4a11 1e-014
Cngan4a7 TDnga13 TDn4a13 1e-014
Cngan4a8 TDnga15 TDn4a15 1e-014
Cngan4a9 TDnga17 TDn4a17 1e-014
Cngan4a10 TDnga19 TDn4a19 1e-014
Cngan4a11 TDnga21 TDn4a21 1e-014
Cngan4a12 TDnga23 TDn4a23 1e-014
Cngan4a13 TDnga25 TDn4a25 1e-014
Cngan4a14 TDnga27 TDn4a27 1e-014
Cngan4a15 TDnga29 TDn4a29 1e-014
Cngan4a16 TDnga31 TDn4a31 1e-014
Cngan4a17 TDnga33 TDn4a33 6e-015
Cngan5a1 TDnga1 TDn5a1 6e-015
Cngan5a2 TDnga3 TDn5a3 1e-014
Cngan5a3 TDnga5 TDn5a5 1e-014
Cngan5a4 TDnga7 TDn5a7 1e-014
Cngan5a5 TDnga9 TDn5a9 1e-014
Cngan5a6 TDnga11 TDn5a11 1e-014
Cngan5a7 TDnga13 TDn5a13 1e-014
Cngan5a8 TDnga15 TDn5a15 1e-014
Cngan5a9 TDnga17 TDn5a17 1e-014
Cngan5a10 TDnga19 TDn5a19 1e-014
Cngan5a11 TDnga21 TDn5a21 1e-014
Cngan5a12 TDnga23 TDn5a23 1e-014
Cngan5a13 TDnga25 TDn5a25 1e-014
Cngan5a14 TDnga27 TDn5a27 1e-014
Cngan5a15 TDnga29 TDn5a29 1e-014
Cngan5a16 TDnga31 TDn5a31 1e-014
Cngan5a17 TDnga33 TDn5a33 6e-015
Cngan6a1 TDnga1 TDn6a1 6e-015
Cngan6a2 TDnga3 TDn6a3 1e-014
Cngan6a3 TDnga5 TDn6a5 1e-014
Cngan6a4 TDnga7 TDn6a7 1e-014
Cngan6a5 TDnga9 TDn6a9 1e-014
Cngan6a6 TDnga11 TDn6a11 1e-014
Cngan6a7 TDnga13 TDn6a13 1e-014
Cngan6a8 TDnga15 TDn6a15 1e-014
Cngan6a9 TDnga17 TDn6a17 1e-014
Cngan6a10 TDnga19 TDn6a19 1e-014
Cngan6a11 TDnga21 TDn6a21 1e-014
Cngan6a12 TDnga23 TDn6a23 1e-014
Cngan6a13 TDnga25 TDn6a25 1e-014
Cngan6a14 TDnga27 TDn6a27 1e-014
Cngan6a15 TDnga29 TDn6a29 1e-014
Cngan6a16 TDnga31 TDn6a31 1e-014
Cngan6a17 TDnga33 TDn6a33 6e-015
Cngan7a1 TDnga1 TDn7a1 5.734420e-015
Cngan7a2 TDnga3 TDn7a3 1e-014
Cngan7a3 TDnga5 TDn7a5 1e-014
Cngan7a4 TDnga7 TDn7a7 1e-014
Cngan7a5 TDnga9 TDn7a9 1e-014
Cngan7a6 TDnga11 TDn7a11 1e-014
Cngan7a7 TDnga13 TDn7a13 1e-014
Cngan7a8 TDnga15 TDn7a15 1e-014
Cngan7a9 TDnga17 TDn7a17 1e-014
Cngan7a10 TDnga19 TDn7a19 1e-014
Cngan7a11 TDnga21 TDn7a21 1e-014
Cngan7a12 TDnga23 TDn7a23 1e-014
Cngan7a13 TDnga25 TDn7a25 1e-014
Cngan7a14 TDnga27 TDn7a27 1e-014
Cngan7a15 TDnga29 TDn7a29 1e-014
Cngan7a16 TDnga31 TDn7a31 1e-014
Cngan7a17 TDnga33 TDn7a33 5.734420e-015
Cngan8a1 TDnga1 TDn8a1 5.773050e-015
Cngan8a2 TDnga3 TDn8a3 1e-014
Cngan8a3 TDnga5 TDn8a5 1e-014
Cngan8a4 TDnga7 TDn8a7 1e-014
Cngan8a5 TDnga9 TDn8a9 1e-014
Cngan8a6 TDnga11 TDn8a11 1e-014
Cngan8a7 TDnga13 TDn8a13 1e-014
Cngan8a8 TDnga15 TDn8a15 1e-014
Cngan8a9 TDnga17 TDn8a17 1e-014
Cngan8a10 TDnga19 TDn8a19 1e-014
Cngan8a11 TDnga21 TDn8a21 1e-014
Cngan8a12 TDnga23 TDn8a23 1e-014
Cngan8a13 TDnga25 TDn8a25 1e-014
Cngan8a14 TDnga27 TDn8a27 1e-014
Cngan8a15 TDnga29 TDn8a29 1e-014
Cngan8a16 TDnga31 TDn8a31 1e-014
Cngan8a17 TDnga33 TDn8a33 5.773050e-015
Cngan9a1 TDnga1 TDn9a1 6.592280e-015
Cngan9a2 TDnga3 TDn9a3 1e-014
Cngan9a3 TDnga5 TDn9a5 1e-014
Cngan9a4 TDnga7 TDn9a7 1e-014
Cngan9a5 TDnga9 TDn9a9 1e-014
Cngan9a6 TDnga11 TDn9a11 1e-014
Cngan9a7 TDnga13 TDn9a13 1e-014
Cngan9a8 TDnga15 TDn9a15 1e-014
Cngan9a9 TDnga17 TDn9a17 1e-014
Cngan9a10 TDnga19 TDn9a19 1e-014
Cngan9a11 TDnga21 TDn9a21 1e-014
Cngan9a12 TDnga23 TDn9a23 1e-014
Cngan9a13 TDnga25 TDn9a25 1e-014
Cngan9a14 TDnga27 TDn9a27 1e-014
Cngan9a15 TDnga29 TDn9a29 1e-014
Cngan9a16 TDnga31 TDn9a31 1e-014
Cngan9a17 TDnga33 TDn9a33 6.592280e-015
Cngan10a1 TDnga1 TDn10a1 2e-014
Cngan10a2 TDnga3 TDn10a3 1e-014
Cngan10a3 TDnga5 TDn10a5 1e-014
Cngan10a4 TDnga7 TDn10a7 1e-014
Cngan10a5 TDnga9 TDn10a9 1e-014
Cngan10a6 TDnga11 TDn10a11 1e-014
Cngan10a7 TDnga13 TDn10a13 1e-014
Cngan10a8 TDnga15 TDn10a15 1e-014
Cngan10a9 TDnga17 TDn10a17 1e-014
Cngan10a10 TDnga19 TDn10a19 1e-014
Cngan10a11 TDnga21 TDn10a21 1e-014
Cngan10a12 TDnga23 TDn10a23 1e-014
Cngan10a13 TDnga25 TDn10a25 1e-014
Cngan10a14 TDnga27 TDn10a27 1e-014
Cngan10a15 TDnga29 TDn10a29 1e-014
Cngan10a16 TDnga31 TDn10a31 1e-014
Cngan10a17 TDnga33 TDn10a33 2e-014
Cngan11a1 TDnga1 TDn11a1 2e-014
Cngan11a2 TDnga3 TDn11a3 1e-014
Cngan11a3 TDnga5 TDn11a5 1e-014
Cngan11a4 TDnga7 TDn11a7 1e-014
Cngan11a5 TDnga9 TDn11a9 1e-014
Cngan11a6 TDnga11 TDn11a11 1e-014
Cngan11a7 TDnga13 TDn11a13 1e-014
Cngan11a8 TDnga15 TDn11a15 1e-014
Cngan11a9 TDnga17 TDn11a17 1e-014
Cngan11a10 TDnga19 TDn11a19 1e-014
Cngan11a11 TDnga21 TDn11a21 1e-014
Cngan11a12 TDnga23 TDn11a23 1e-014
Cngan11a13 TDnga25 TDn11a25 1e-014
Cngan11a14 TDnga27 TDn11a27 1e-014
Cngan11a15 TDnga29 TDn11a29 1e-014
Cngan11a16 TDnga31 TDn11a31 1e-014
Cngan11a17 TDnga33 TDn11a33 2e-014
Cngan12a1 TDnga1 TDn12a1 2e-014
Cngan12a2 TDnga3 TDn12a3 1e-014
Cngan12a3 TDnga5 TDn12a5 1e-014
Cngan12a4 TDnga7 TDn12a7 1e-014
Cngan12a5 TDnga9 TDn12a9 1e-014
Cngan12a6 TDnga11 TDn12a11 1e-014
Cngan12a7 TDnga13 TDn12a13 1e-014
Cngan12a8 TDnga15 TDn12a15 1e-014
Cngan12a9 TDnga17 TDn12a17 1e-014
Cngan12a10 TDnga19 TDn12a19 1e-014
Cngan12a11 TDnga21 TDn12a21 1e-014
Cngan12a12 TDnga23 TDn12a23 1e-014
Cngan12a13 TDnga25 TDn12a25 1e-014
Cngan12a14 TDnga27 TDn12a27 1e-014
Cngan12a15 TDnga29 TDn12a29 1e-014
Cngan12a16 TDnga31 TDn12a31 1e-014
Cngan12a17 TDnga33 TDn12a33 2e-014
Cnganva1 TDnga1 TDnva1 2e-014
Cnganva2 TDnga3 TDnva3 1e-014
Cnganva3 TDnga5 TDnva5 1e-014
Cnganva4 TDnga7 TDnva7 1e-014
Cnganva5 TDnga9 TDnva9 1e-014
Cnganva6 TDnga11 TDnva11 1e-014
Cnganva7 TDnga13 TDnva13 1e-014
Cnganva8 TDnga15 TDnva15 1e-014
Cnganva9 TDnga17 TDnva17 1e-014
Cnganva10 TDnga19 TDnva19 1e-014
Cnganva11 TDnga21 TDnva21 1e-014
Cnganva12 TDnga23 TDnva23 1e-014
Cnganva13 TDnga25 TDnva25 1e-014
Cnganva14 TDnga27 TDnva27 1e-014
Cnganva15 TDnga29 TDnva29 1e-014
Cnganva16 TDnga31 TDnva31 1e-014
Cnganva17 TDnga33 TDnva33 2e-014
Cn1an2a1 TDn1a1 TDn2a1 1.586220e-014
Cn1an2a2 TDn1a3 TDn2a3 3e-014
Cn1an2a3 TDn1a5 TDn2a5 3e-014
Cn1an2a4 TDn1a7 TDn2a7 3e-014
Cn1an2a5 TDn1a9 TDn2a9 3e-014
Cn1an2a6 TDn1a11 TDn2a11 3e-014
Cn1an2a7 TDn1a13 TDn2a13 3e-014
Cn1an2a8 TDn1a15 TDn2a15 3e-014
Cn1an2a9 TDn1a17 TDn2a17 3e-014
Cn1an2a10 TDn1a19 TDn2a19 3e-014
Cn1an2a11 TDn1a21 TDn2a21 3e-014
Cn1an2a12 TDn1a23 TDn2a23 3e-014
Cn1an2a13 TDn1a25 TDn2a25 3e-014
Cn1an2a14 TDn1a27 TDn2a27 3e-014
Cn1an2a15 TDn1a29 TDn2a29 3e-014
Cn1an2a16 TDn1a31 TDn2a31 3e-014
Cn1an2a17 TDn1a33 TDn2a33 1.586220e-014
Cn1an3a1 TDn1a1 TDn3a1 5.674250e-015
Cn1an3a2 TDn1a3 TDn3a3 1e-014
Cn1an3a3 TDn1a5 TDn3a5 1e-014
Cn1an3a4 TDn1a7 TDn3a7 1e-014
Cn1an3a5 TDn1a9 TDn3a9 1e-014
Cn1an3a6 TDn1a11 TDn3a11 1e-014
Cn1an3a7 TDn1a13 TDn3a13 1e-014
Cn1an3a8 TDn1a15 TDn3a15 1e-014
Cn1an3a9 TDn1a17 TDn3a17 1e-014
Cn1an3a10 TDn1a19 TDn3a19 1e-014
Cn1an3a11 TDn1a21 TDn3a21 1e-014
Cn1an3a12 TDn1a23 TDn3a23 1e-014
Cn1an3a13 TDn1a25 TDn3a25 1e-014
Cn1an3a14 TDn1a27 TDn3a27 1e-014
Cn1an3a15 TDn1a29 TDn3a29 1e-014
Cn1an3a16 TDn1a31 TDn3a31 1e-014
Cn1an3a17 TDn1a33 TDn3a33 5.674250e-015
Cn1an4a1 TDn1a1 TDn4a1 5.219520e-015
Cn1an4a2 TDn1a3 TDn4a3 1e-014
Cn1an4a3 TDn1a5 TDn4a5 1e-014
Cn1an4a4 TDn1a7 TDn4a7 1e-014
Cn1an4a5 TDn1a9 TDn4a9 1e-014
Cn1an4a6 TDn1a11 TDn4a11 1e-014
Cn1an4a7 TDn1a13 TDn4a13 1e-014
Cn1an4a8 TDn1a15 TDn4a15 1e-014
Cn1an4a9 TDn1a17 TDn4a17 1e-014
Cn1an4a10 TDn1a19 TDn4a19 1e-014
Cn1an4a11 TDn1a21 TDn4a21 1e-014
Cn1an4a12 TDn1a23 TDn4a23 1e-014
Cn1an4a13 TDn1a25 TDn4a25 1e-014
Cn1an4a14 TDn1a27 TDn4a27 1e-014
Cn1an4a15 TDn1a29 TDn4a29 1e-014
Cn1an4a16 TDn1a31 TDn4a31 1e-014
Cn1an4a17 TDn1a33 TDn4a33 5.219520e-015
Cn1an5a1 TDn1a1 TDn5a1 5.062210e-015
Cn1an5a2 TDn1a3 TDn5a3 1e-014
Cn1an5a3 TDn1a5 TDn5a5 1e-014
Cn1an5a4 TDn1a7 TDn5a7 1e-014
Cn1an5a5 TDn1a9 TDn5a9 1e-014
Cn1an5a6 TDn1a11 TDn5a11 1e-014
Cn1an5a7 TDn1a13 TDn5a13 1e-014
Cn1an5a8 TDn1a15 TDn5a15 1e-014
Cn1an5a9 TDn1a17 TDn5a17 1e-014
Cn1an5a10 TDn1a19 TDn5a19 1e-014
Cn1an5a11 TDn1a21 TDn5a21 1e-014
Cn1an5a12 TDn1a23 TDn5a23 1e-014
Cn1an5a13 TDn1a25 TDn5a25 1e-014
Cn1an5a14 TDn1a27 TDn5a27 1e-014
Cn1an5a15 TDn1a29 TDn5a29 1e-014
Cn1an5a16 TDn1a31 TDn5a31 1e-014
Cn1an5a17 TDn1a33 TDn5a33 5.062210e-015
Cn1an6a1 TDn1a1 TDn6a1 5.003840e-015
Cn1an6a2 TDn1a3 TDn6a3 1e-014
Cn1an6a3 TDn1a5 TDn6a5 1e-014
Cn1an6a4 TDn1a7 TDn6a7 1e-014
Cn1an6a5 TDn1a9 TDn6a9 1e-014
Cn1an6a6 TDn1a11 TDn6a11 1e-014
Cn1an6a7 TDn1a13 TDn6a13 1e-014
Cn1an6a8 TDn1a15 TDn6a15 1e-014
Cn1an6a9 TDn1a17 TDn6a17 1e-014
Cn1an6a10 TDn1a19 TDn6a19 1e-014
Cn1an6a11 TDn1a21 TDn6a21 1e-014
Cn1an6a12 TDn1a23 TDn6a23 1e-014
Cn1an6a13 TDn1a25 TDn6a25 1e-014
Cn1an6a14 TDn1a27 TDn6a27 1e-014
Cn1an6a15 TDn1a29 TDn6a29 1e-014
Cn1an6a16 TDn1a31 TDn6a31 1e-014
Cn1an6a17 TDn1a33 TDn6a33 5.003840e-015
Cn1an7a1 TDn1a1 TDn7a1 4.990870e-015
Cn1an7a2 TDn1a3 TDn7a3 1e-014
Cn1an7a3 TDn1a5 TDn7a5 1e-014
Cn1an7a4 TDn1a7 TDn7a7 1e-014
Cn1an7a5 TDn1a9 TDn7a9 1e-014
Cn1an7a6 TDn1a11 TDn7a11 1e-014
Cn1an7a7 TDn1a13 TDn7a13 1e-014
Cn1an7a8 TDn1a15 TDn7a15 1e-014
Cn1an7a9 TDn1a17 TDn7a17 1e-014
Cn1an7a10 TDn1a19 TDn7a19 1e-014
Cn1an7a11 TDn1a21 TDn7a21 1e-014
Cn1an7a12 TDn1a23 TDn7a23 1e-014
Cn1an7a13 TDn1a25 TDn7a25 1e-014
Cn1an7a14 TDn1a27 TDn7a27 1e-014
Cn1an7a15 TDn1a29 TDn7a29 1e-014
Cn1an7a16 TDn1a31 TDn7a31 1e-014
Cn1an7a17 TDn1a33 TDn7a33 4.990870e-015
Cn1an8a1 TDn1a1 TDn8a1 5.026740e-015
Cn1an8a2 TDn1a3 TDn8a3 1e-014
Cn1an8a3 TDn1a5 TDn8a5 1e-014
Cn1an8a4 TDn1a7 TDn8a7 1e-014
Cn1an8a5 TDn1a9 TDn8a9 1e-014
Cn1an8a6 TDn1a11 TDn8a11 1e-014
Cn1an8a7 TDn1a13 TDn8a13 1e-014
Cn1an8a8 TDn1a15 TDn8a15 1e-014
Cn1an8a9 TDn1a17 TDn8a17 1e-014
Cn1an8a10 TDn1a19 TDn8a19 1e-014
Cn1an8a11 TDn1a21 TDn8a21 1e-014
Cn1an8a12 TDn1a23 TDn8a23 1e-014
Cn1an8a13 TDn1a25 TDn8a25 1e-014
Cn1an8a14 TDn1a27 TDn8a27 1e-014
Cn1an8a15 TDn1a29 TDn8a29 1e-014
Cn1an8a16 TDn1a31 TDn8a31 1e-014
Cn1an8a17 TDn1a33 TDn8a33 5.026740e-015
Cn1an9a1 TDn1a1 TDn9a1 5.751040e-015
Cn1an9a2 TDn1a3 TDn9a3 1e-014
Cn1an9a3 TDn1a5 TDn9a5 1e-014
Cn1an9a4 TDn1a7 TDn9a7 1e-014
Cn1an9a5 TDn1a9 TDn9a9 1e-014
Cn1an9a6 TDn1a11 TDn9a11 1e-014
Cn1an9a7 TDn1a13 TDn9a13 1e-014
Cn1an9a8 TDn1a15 TDn9a15 1e-014
Cn1an9a9 TDn1a17 TDn9a17 1e-014
Cn1an9a10 TDn1a19 TDn9a19 1e-014
Cn1an9a11 TDn1a21 TDn9a21 1e-014
Cn1an9a12 TDn1a23 TDn9a23 1e-014
Cn1an9a13 TDn1a25 TDn9a25 1e-014
Cn1an9a14 TDn1a27 TDn9a27 1e-014
Cn1an9a15 TDn1a29 TDn9a29 1e-014
Cn1an9a16 TDn1a31 TDn9a31 1e-014
Cn1an9a17 TDn1a33 TDn9a33 5.751040e-015
Cn1an10a1 TDn1a1 TDn10a1 2e-014
Cn1an10a2 TDn1a3 TDn10a3 1e-014
Cn1an10a3 TDn1a5 TDn10a5 1e-014
Cn1an10a4 TDn1a7 TDn10a7 1e-014
Cn1an10a5 TDn1a9 TDn10a9 1e-014
Cn1an10a6 TDn1a11 TDn10a11 1e-014
Cn1an10a7 TDn1a13 TDn10a13 1e-014
Cn1an10a8 TDn1a15 TDn10a15 1e-014
Cn1an10a9 TDn1a17 TDn10a17 1e-014
Cn1an10a10 TDn1a19 TDn10a19 1e-014
Cn1an10a11 TDn1a21 TDn10a21 1e-014
Cn1an10a12 TDn1a23 TDn10a23 1e-014
Cn1an10a13 TDn1a25 TDn10a25 1e-014
Cn1an10a14 TDn1a27 TDn10a27 1e-014
Cn1an10a15 TDn1a29 TDn10a29 1e-014
Cn1an10a16 TDn1a31 TDn10a31 1e-014
Cn1an10a17 TDn1a33 TDn10a33 2e-014
Cn1an11a1 TDn1a1 TDn11a1 2e-014
Cn1an11a2 TDn1a3 TDn11a3 1e-014
Cn1an11a3 TDn1a5 TDn11a5 1e-014
Cn1an11a4 TDn1a7 TDn11a7 1e-014
Cn1an11a5 TDn1a9 TDn11a9 1e-014
Cn1an11a6 TDn1a11 TDn11a11 1e-014
Cn1an11a7 TDn1a13 TDn11a13 1e-014
Cn1an11a8 TDn1a15 TDn11a15 1e-014
Cn1an11a9 TDn1a17 TDn11a17 1e-014
Cn1an11a10 TDn1a19 TDn11a19 1e-014
Cn1an11a11 TDn1a21 TDn11a21 1e-014
Cn1an11a12 TDn1a23 TDn11a23 1e-014
Cn1an11a13 TDn1a25 TDn11a25 1e-014
Cn1an11a14 TDn1a27 TDn11a27 1e-014
Cn1an11a15 TDn1a29 TDn11a29 1e-014
Cn1an11a16 TDn1a31 TDn11a31 1e-014
Cn1an11a17 TDn1a33 TDn11a33 2e-014
Cn1an12a1 TDn1a1 TDn12a1 2e-014
Cn1an12a2 TDn1a3 TDn12a3 1e-014
Cn1an12a3 TDn1a5 TDn12a5 1e-014
Cn1an12a4 TDn1a7 TDn12a7 1e-014
Cn1an12a5 TDn1a9 TDn12a9 1e-014
Cn1an12a6 TDn1a11 TDn12a11 1e-014
Cn1an12a7 TDn1a13 TDn12a13 1e-014
Cn1an12a8 TDn1a15 TDn12a15 1e-014
Cn1an12a9 TDn1a17 TDn12a17 1e-014
Cn1an12a10 TDn1a19 TDn12a19 1e-014
Cn1an12a11 TDn1a21 TDn12a21 1e-014
Cn1an12a12 TDn1a23 TDn12a23 1e-014
Cn1an12a13 TDn1a25 TDn12a25 1e-014
Cn1an12a14 TDn1a27 TDn12a27 1e-014
Cn1an12a15 TDn1a29 TDn12a29 1e-014
Cn1an12a16 TDn1a31 TDn12a31 1e-014
Cn1an12a17 TDn1a33 TDn12a33 2e-014
Cn1anva1 TDn1a1 TDnva1 2e-014
Cn1anva2 TDn1a3 TDnva3 2e-014
Cn1anva3 TDn1a5 TDnva5 2e-014
Cn1anva4 TDn1a7 TDnva7 2e-014
Cn1anva5 TDn1a9 TDnva9 2e-014
Cn1anva6 TDn1a11 TDnva11 2e-014
Cn1anva7 TDn1a13 TDnva13 2e-014
Cn1anva8 TDn1a15 TDnva15 2e-014
Cn1anva9 TDn1a17 TDnva17 2e-014
Cn1anva10 TDn1a19 TDnva19 2e-014
Cn1anva11 TDn1a21 TDnva21 2e-014
Cn1anva12 TDn1a23 TDnva23 2e-014
Cn1anva13 TDn1a25 TDnva25 2e-014
Cn1anva14 TDn1a27 TDnva27 2e-014
Cn1anva15 TDn1a29 TDnva29 2e-014
Cn1anva16 TDn1a31 TDnva31 2e-014
Cn1anva17 TDn1a33 TDnva33 2e-014
Cn2an3a1 TDn2a1 TDn3a1 1.576950e-014
Cn2an3a2 TDn2a3 TDn3a3 3.153910e-014
Cn2an3a3 TDn2a5 TDn3a5 3.153910e-014
Cn2an3a4 TDn2a7 TDn3a7 3.153910e-014
Cn2an3a5 TDn2a9 TDn3a9 3.153910e-014
Cn2an3a6 TDn2a11 TDn3a11 3.153910e-014
Cn2an3a7 TDn2a13 TDn3a13 3.153910e-014
Cn2an3a8 TDn2a15 TDn3a15 3.153910e-014
Cn2an3a9 TDn2a17 TDn3a17 3.153910e-014
Cn2an3a10 TDn2a19 TDn3a19 3.153910e-014
Cn2an3a11 TDn2a21 TDn3a21 3.153910e-014
Cn2an3a12 TDn2a23 TDn3a23 3.153910e-014
Cn2an3a13 TDn2a25 TDn3a25 3.153910e-014
Cn2an3a14 TDn2a27 TDn3a27 3.153910e-014
Cn2an3a15 TDn2a29 TDn3a29 3.153910e-014
Cn2an3a16 TDn2a31 TDn3a31 3.153910e-014
Cn2an3a17 TDn2a33 TDn3a33 1.576950e-014
Cn2an4a1 TDn2a1 TDn4a1 5.623050e-015
Cn2an4a2 TDn2a3 TDn4a3 1e-014
Cn2an4a3 TDn2a5 TDn4a5 1e-014
Cn2an4a4 TDn2a7 TDn4a7 1e-014
Cn2an4a5 TDn2a9 TDn4a9 1e-014
Cn2an4a6 TDn2a11 TDn4a11 1e-014
Cn2an4a7 TDn2a13 TDn4a13 1e-014
Cn2an4a8 TDn2a15 TDn4a15 1e-014
Cn2an4a9 TDn2a17 TDn4a17 1e-014
Cn2an4a10 TDn2a19 TDn4a19 1e-014
Cn2an4a11 TDn2a21 TDn4a21 1e-014
Cn2an4a12 TDn2a23 TDn4a23 1e-014
Cn2an4a13 TDn2a25 TDn4a25 1e-014
Cn2an4a14 TDn2a27 TDn4a27 1e-014
Cn2an4a15 TDn2a29 TDn4a29 1e-014
Cn2an4a16 TDn2a31 TDn4a31 1e-014
Cn2an4a17 TDn2a33 TDn4a33 5.623050e-015
Cn2an5a1 TDn2a1 TDn5a1 5.149670e-015
Cn2an5a2 TDn2a3 TDn5a3 1e-014
Cn2an5a3 TDn2a5 TDn5a5 1e-014
Cn2an5a4 TDn2a7 TDn5a7 1e-014
Cn2an5a5 TDn2a9 TDn5a9 1e-014
Cn2an5a6 TDn2a11 TDn5a11 1e-014
Cn2an5a7 TDn2a13 TDn5a13 1e-014
Cn2an5a8 TDn2a15 TDn5a15 1e-014
Cn2an5a9 TDn2a17 TDn5a17 1e-014
Cn2an5a10 TDn2a19 TDn5a19 1e-014
Cn2an5a11 TDn2a21 TDn5a21 1e-014
Cn2an5a12 TDn2a23 TDn5a23 1e-014
Cn2an5a13 TDn2a25 TDn5a25 1e-014
Cn2an5a14 TDn2a27 TDn5a27 1e-014
Cn2an5a15 TDn2a29 TDn5a29 1e-014
Cn2an5a16 TDn2a31 TDn5a31 1e-014
Cn2an5a17 TDn2a33 TDn5a33 5.149670e-015
Cn2an6a1 TDn2a1 TDn6a1 5.011480e-015
Cn2an6a2 TDn2a3 TDn6a3 1e-014
Cn2an6a3 TDn2a5 TDn6a5 1e-014
Cn2an6a4 TDn2a7 TDn6a7 1e-014
Cn2an6a5 TDn2a9 TDn6a9 1e-014
Cn2an6a6 TDn2a11 TDn6a11 1e-014
Cn2an6a7 TDn2a13 TDn6a13 1e-014
Cn2an6a8 TDn2a15 TDn6a15 1e-014
Cn2an6a9 TDn2a17 TDn6a17 1e-014
Cn2an6a10 TDn2a19 TDn6a19 1e-014
Cn2an6a11 TDn2a21 TDn6a21 1e-014
Cn2an6a12 TDn2a23 TDn6a23 1e-014
Cn2an6a13 TDn2a25 TDn6a25 1e-014
Cn2an6a14 TDn2a27 TDn6a27 1e-014
Cn2an6a15 TDn2a29 TDn6a29 1e-014
Cn2an6a16 TDn2a31 TDn6a31 1e-014
Cn2an6a17 TDn2a33 TDn6a33 5.011480e-015
Cn2an7a1 TDn2a1 TDn7a1 4.968610e-015
Cn2an7a2 TDn2a3 TDn7a3 1e-014
Cn2an7a3 TDn2a5 TDn7a5 1e-014
Cn2an7a4 TDn2a7 TDn7a7 1e-014
Cn2an7a5 TDn2a9 TDn7a9 1e-014
Cn2an7a6 TDn2a11 TDn7a11 1e-014
Cn2an7a7 TDn2a13 TDn7a13 1e-014
Cn2an7a8 TDn2a15 TDn7a15 1e-014
Cn2an7a9 TDn2a17 TDn7a17 1e-014
Cn2an7a10 TDn2a19 TDn7a19 1e-014
Cn2an7a11 TDn2a21 TDn7a21 1e-014
Cn2an7a12 TDn2a23 TDn7a23 1e-014
Cn2an7a13 TDn2a25 TDn7a25 1e-014
Cn2an7a14 TDn2a27 TDn7a27 1e-014
Cn2an7a15 TDn2a29 TDn7a29 1e-014
Cn2an7a16 TDn2a31 TDn7a31 1e-014
Cn2an7a17 TDn2a33 TDn7a33 4.968610e-015
Cn2an8a1 TDn2a1 TDn8a1 4.990350e-015
Cn2an8a2 TDn2a3 TDn8a3 1e-014
Cn2an8a3 TDn2a5 TDn8a5 1e-014
Cn2an8a4 TDn2a7 TDn8a7 1e-014
Cn2an8a5 TDn2a9 TDn8a9 1e-014
Cn2an8a6 TDn2a11 TDn8a11 1e-014
Cn2an8a7 TDn2a13 TDn8a13 1e-014
Cn2an8a8 TDn2a15 TDn8a15 1e-014
Cn2an8a9 TDn2a17 TDn8a17 1e-014
Cn2an8a10 TDn2a19 TDn8a19 1e-014
Cn2an8a11 TDn2a21 TDn8a21 1e-014
Cn2an8a12 TDn2a23 TDn8a23 1e-014
Cn2an8a13 TDn2a25 TDn8a25 1e-014
Cn2an8a14 TDn2a27 TDn8a27 1e-014
Cn2an8a15 TDn2a29 TDn8a29 1e-014
Cn2an8a16 TDn2a31 TDn8a31 1e-014
Cn2an8a17 TDn2a33 TDn8a33 4.990350e-015
Cn2an9a1 TDn2a1 TDn9a1 5.701980e-015
Cn2an9a2 TDn2a3 TDn9a3 1e-014
Cn2an9a3 TDn2a5 TDn9a5 1e-014
Cn2an9a4 TDn2a7 TDn9a7 1e-014
Cn2an9a5 TDn2a9 TDn9a9 1e-014
Cn2an9a6 TDn2a11 TDn9a11 1e-014
Cn2an9a7 TDn2a13 TDn9a13 1e-014
Cn2an9a8 TDn2a15 TDn9a15 1e-014
Cn2an9a9 TDn2a17 TDn9a17 1e-014
Cn2an9a10 TDn2a19 TDn9a19 1e-014
Cn2an9a11 TDn2a21 TDn9a21 1e-014
Cn2an9a12 TDn2a23 TDn9a23 1e-014
Cn2an9a13 TDn2a25 TDn9a25 1e-014
Cn2an9a14 TDn2a27 TDn9a27 1e-014
Cn2an9a15 TDn2a29 TDn9a29 1e-014
Cn2an9a16 TDn2a31 TDn9a31 1e-014
Cn2an9a17 TDn2a33 TDn9a33 5.701980e-015
Cn2an10a1 TDn2a1 TDn10a1 2e-014
Cn2an10a2 TDn2a3 TDn10a3 1e-014
Cn2an10a3 TDn2a5 TDn10a5 1e-014
Cn2an10a4 TDn2a7 TDn10a7 1e-014
Cn2an10a5 TDn2a9 TDn10a9 1e-014
Cn2an10a6 TDn2a11 TDn10a11 1e-014
Cn2an10a7 TDn2a13 TDn10a13 1e-014
Cn2an10a8 TDn2a15 TDn10a15 1e-014
Cn2an10a9 TDn2a17 TDn10a17 1e-014
Cn2an10a10 TDn2a19 TDn10a19 1e-014
Cn2an10a11 TDn2a21 TDn10a21 1e-014
Cn2an10a12 TDn2a23 TDn10a23 1e-014
Cn2an10a13 TDn2a25 TDn10a25 1e-014
Cn2an10a14 TDn2a27 TDn10a27 1e-014
Cn2an10a15 TDn2a29 TDn10a29 1e-014
Cn2an10a16 TDn2a31 TDn10a31 1e-014
Cn2an10a17 TDn2a33 TDn10a33 2e-014
Cn2an11a1 TDn2a1 TDn11a1 2e-014
Cn2an11a2 TDn2a3 TDn11a3 1e-014
Cn2an11a3 TDn2a5 TDn11a5 1e-014
Cn2an11a4 TDn2a7 TDn11a7 1e-014
Cn2an11a5 TDn2a9 TDn11a9 1e-014
Cn2an11a6 TDn2a11 TDn11a11 1e-014
Cn2an11a7 TDn2a13 TDn11a13 1e-014
Cn2an11a8 TDn2a15 TDn11a15 1e-014
Cn2an11a9 TDn2a17 TDn11a17 1e-014
Cn2an11a10 TDn2a19 TDn11a19 1e-014
Cn2an11a11 TDn2a21 TDn11a21 1e-014
Cn2an11a12 TDn2a23 TDn11a23 1e-014
Cn2an11a13 TDn2a25 TDn11a25 1e-014
Cn2an11a14 TDn2a27 TDn11a27 1e-014
Cn2an11a15 TDn2a29 TDn11a29 1e-014
Cn2an11a16 TDn2a31 TDn11a31 1e-014
Cn2an11a17 TDn2a33 TDn11a33 2e-014
Cn2an12a1 TDn2a1 TDn12a1 2e-014
Cn2an12a2 TDn2a3 TDn12a3 1e-014
Cn2an12a3 TDn2a5 TDn12a5 1e-014
Cn2an12a4 TDn2a7 TDn12a7 1e-014
Cn2an12a5 TDn2a9 TDn12a9 1e-014
Cn2an12a6 TDn2a11 TDn12a11 1e-014
Cn2an12a7 TDn2a13 TDn12a13 1e-014
Cn2an12a8 TDn2a15 TDn12a15 1e-014
Cn2an12a9 TDn2a17 TDn12a17 1e-014
Cn2an12a10 TDn2a19 TDn12a19 1e-014
Cn2an12a11 TDn2a21 TDn12a21 1e-014
Cn2an12a12 TDn2a23 TDn12a23 1e-014
Cn2an12a13 TDn2a25 TDn12a25 1e-014
Cn2an12a14 TDn2a27 TDn12a27 1e-014
Cn2an12a15 TDn2a29 TDn12a29 1e-014
Cn2an12a16 TDn2a31 TDn12a31 1e-014
Cn2an12a17 TDn2a33 TDn12a33 2e-014
Cn2anva1 TDn2a1 TDnva1 2e-014
Cn2anva2 TDn2a3 TDnva3 2e-014
Cn2anva3 TDn2a5 TDnva5 2e-014
Cn2anva4 TDn2a7 TDnva7 2e-014
Cn2anva5 TDn2a9 TDnva9 2e-014
Cn2anva6 TDn2a11 TDnva11 2e-014
Cn2anva7 TDn2a13 TDnva13 2e-014
Cn2anva8 TDn2a15 TDnva15 2e-014
Cn2anva9 TDn2a17 TDnva17 2e-014
Cn2anva10 TDn2a19 TDnva19 2e-014
Cn2anva11 TDn2a21 TDnva21 2e-014
Cn2anva12 TDn2a23 TDnva23 2e-014
Cn2anva13 TDn2a25 TDnva25 2e-014
Cn2anva14 TDn2a27 TDnva27 2e-014
Cn2anva15 TDn2a29 TDnva29 2e-014
Cn2anva16 TDn2a31 TDnva31 2e-014
Cn2anva17 TDn2a33 TDnva33 2e-014
Cn3an4a1 TDn3a1 TDn4a1 1.575450e-014
Cn3an4a2 TDn3a3 TDn4a3 3e-014
Cn3an4a3 TDn3a5 TDn4a5 3e-014
Cn3an4a4 TDn3a7 TDn4a7 3e-014
Cn3an4a5 TDn3a9 TDn4a9 3e-014
Cn3an4a6 TDn3a11 TDn4a11 3e-014
Cn3an4a7 TDn3a13 TDn4a13 3e-014
Cn3an4a8 TDn3a15 TDn4a15 3e-014
Cn3an4a9 TDn3a17 TDn4a17 3e-014
Cn3an4a10 TDn3a19 TDn4a19 3e-014
Cn3an4a11 TDn3a21 TDn4a21 3e-014
Cn3an4a12 TDn3a23 TDn4a23 3e-014
Cn3an4a13 TDn3a25 TDn4a25 3e-014
Cn3an4a14 TDn3a27 TDn4a27 3e-014
Cn3an4a15 TDn3a29 TDn4a29 3e-014
Cn3an4a16 TDn3a31 TDn4a31 3e-014
Cn3an4a17 TDn3a33 TDn4a33 1.575450e-014
Cn3an5a1 TDn3a1 TDn5a1 5.588630e-015
Cn3an5a2 TDn3a3 TDn5a3 1e-014
Cn3an5a3 TDn3a5 TDn5a5 1e-014
Cn3an5a4 TDn3a7 TDn5a7 1e-014
Cn3an5a5 TDn3a9 TDn5a9 1e-014
Cn3an5a6 TDn3a11 TDn5a11 1e-014
Cn3an5a7 TDn3a13 TDn5a13 1e-014
Cn3an5a8 TDn3a15 TDn5a15 1e-014
Cn3an5a9 TDn3a17 TDn5a17 1e-014
Cn3an5a10 TDn3a19 TDn5a19 1e-014
Cn3an5a11 TDn3a21 TDn5a21 1e-014
Cn3an5a12 TDn3a23 TDn5a23 1e-014
Cn3an5a13 TDn3a25 TDn5a25 1e-014
Cn3an5a14 TDn3a27 TDn5a27 1e-014
Cn3an5a15 TDn3a29 TDn5a29 1e-014
Cn3an5a16 TDn3a31 TDn5a31 1e-014
Cn3an5a17 TDn3a33 TDn5a33 5.588630e-015
Cn3an6a1 TDn3a1 TDn6a1 5.135110e-015
Cn3an6a2 TDn3a3 TDn6a3 1e-014
Cn3an6a3 TDn3a5 TDn6a5 1e-014
Cn3an6a4 TDn3a7 TDn6a7 1e-014
Cn3an6a5 TDn3a9 TDn6a9 1e-014
Cn3an6a6 TDn3a11 TDn6a11 1e-014
Cn3an6a7 TDn3a13 TDn6a13 1e-014
Cn3an6a8 TDn3a15 TDn6a15 1e-014
Cn3an6a9 TDn3a17 TDn6a17 1e-014
Cn3an6a10 TDn3a19 TDn6a19 1e-014
Cn3an6a11 TDn3a21 TDn6a21 1e-014
Cn3an6a12 TDn3a23 TDn6a23 1e-014
Cn3an6a13 TDn3a25 TDn6a25 1e-014
Cn3an6a14 TDn3a27 TDn6a27 1e-014
Cn3an6a15 TDn3a29 TDn6a29 1e-014
Cn3an6a16 TDn3a31 TDn6a31 1e-014
Cn3an6a17 TDn3a33 TDn6a33 5.135110e-015
Cn3an7a1 TDn3a1 TDn7a1 5.012180e-015
Cn3an7a2 TDn3a3 TDn7a3 1e-014
Cn3an7a3 TDn3a5 TDn7a5 1e-014
Cn3an7a4 TDn3a7 TDn7a7 1e-014
Cn3an7a5 TDn3a9 TDn7a9 1e-014
Cn3an7a6 TDn3a11 TDn7a11 1e-014
Cn3an7a7 TDn3a13 TDn7a13 1e-014
Cn3an7a8 TDn3a15 TDn7a15 1e-014
Cn3an7a9 TDn3a17 TDn7a17 1e-014
Cn3an7a10 TDn3a19 TDn7a19 1e-014
Cn3an7a11 TDn3a21 TDn7a21 1e-014
Cn3an7a12 TDn3a23 TDn7a23 1e-014
Cn3an7a13 TDn3a25 TDn7a25 1e-014
Cn3an7a14 TDn3a27 TDn7a27 1e-014
Cn3an7a15 TDn3a29 TDn7a29 1e-014
Cn3an7a16 TDn3a31 TDn7a31 1e-014
Cn3an7a17 TDn3a33 TDn7a33 5.012180e-015
Cn3an8a1 TDn3a1 TDn8a1 5.004030e-015
Cn3an8a2 TDn3a3 TDn8a3 1e-014
Cn3an8a3 TDn3a5 TDn8a5 1e-014
Cn3an8a4 TDn3a7 TDn8a7 1e-014
Cn3an8a5 TDn3a9 TDn8a9 1e-014
Cn3an8a6 TDn3a11 TDn8a11 1e-014
Cn3an8a7 TDn3a13 TDn8a13 1e-014
Cn3an8a8 TDn3a15 TDn8a15 1e-014
Cn3an8a9 TDn3a17 TDn8a17 1e-014
Cn3an8a10 TDn3a19 TDn8a19 1e-014
Cn3an8a11 TDn3a21 TDn8a21 1e-014
Cn3an8a12 TDn3a23 TDn8a23 1e-014
Cn3an8a13 TDn3a25 TDn8a25 1e-014
Cn3an8a14 TDn3a27 TDn8a27 1e-014
Cn3an8a15 TDn3a29 TDn8a29 1e-014
Cn3an8a16 TDn3a31 TDn8a31 1e-014
Cn3an8a17 TDn3a33 TDn8a33 5.004030e-015
Cn3an9a1 TDn3a1 TDn9a1 5.703560e-015
Cn3an9a2 TDn3a3 TDn9a3 1e-014
Cn3an9a3 TDn3a5 TDn9a5 1e-014
Cn3an9a4 TDn3a7 TDn9a7 1e-014
Cn3an9a5 TDn3a9 TDn9a9 1e-014
Cn3an9a6 TDn3a11 TDn9a11 1e-014
Cn3an9a7 TDn3a13 TDn9a13 1e-014
Cn3an9a8 TDn3a15 TDn9a15 1e-014
Cn3an9a9 TDn3a17 TDn9a17 1e-014
Cn3an9a10 TDn3a19 TDn9a19 1e-014
Cn3an9a11 TDn3a21 TDn9a21 1e-014
Cn3an9a12 TDn3a23 TDn9a23 1e-014
Cn3an9a13 TDn3a25 TDn9a25 1e-014
Cn3an9a14 TDn3a27 TDn9a27 1e-014
Cn3an9a15 TDn3a29 TDn9a29 1e-014
Cn3an9a16 TDn3a31 TDn9a31 1e-014
Cn3an9a17 TDn3a33 TDn9a33 5.703560e-015
Cn3an10a1 TDn3a1 TDn10a1 2e-014
Cn3an10a2 TDn3a3 TDn10a3 1e-014
Cn3an10a3 TDn3a5 TDn10a5 1e-014
Cn3an10a4 TDn3a7 TDn10a7 1e-014
Cn3an10a5 TDn3a9 TDn10a9 1e-014
Cn3an10a6 TDn3a11 TDn10a11 1e-014
Cn3an10a7 TDn3a13 TDn10a13 1e-014
Cn3an10a8 TDn3a15 TDn10a15 1e-014
Cn3an10a9 TDn3a17 TDn10a17 1e-014
Cn3an10a10 TDn3a19 TDn10a19 1e-014
Cn3an10a11 TDn3a21 TDn10a21 1e-014
Cn3an10a12 TDn3a23 TDn10a23 1e-014
Cn3an10a13 TDn3a25 TDn10a25 1e-014
Cn3an10a14 TDn3a27 TDn10a27 1e-014
Cn3an10a15 TDn3a29 TDn10a29 1e-014
Cn3an10a16 TDn3a31 TDn10a31 1e-014
Cn3an10a17 TDn3a33 TDn10a33 2e-014
Cn3an11a1 TDn3a1 TDn11a1 2e-014
Cn3an11a2 TDn3a3 TDn11a3 1e-014
Cn3an11a3 TDn3a5 TDn11a5 1e-014
Cn3an11a4 TDn3a7 TDn11a7 1e-014
Cn3an11a5 TDn3a9 TDn11a9 1e-014
Cn3an11a6 TDn3a11 TDn11a11 1e-014
Cn3an11a7 TDn3a13 TDn11a13 1e-014
Cn3an11a8 TDn3a15 TDn11a15 1e-014
Cn3an11a9 TDn3a17 TDn11a17 1e-014
Cn3an11a10 TDn3a19 TDn11a19 1e-014
Cn3an11a11 TDn3a21 TDn11a21 1e-014
Cn3an11a12 TDn3a23 TDn11a23 1e-014
Cn3an11a13 TDn3a25 TDn11a25 1e-014
Cn3an11a14 TDn3a27 TDn11a27 1e-014
Cn3an11a15 TDn3a29 TDn11a29 1e-014
Cn3an11a16 TDn3a31 TDn11a31 1e-014
Cn3an11a17 TDn3a33 TDn11a33 2e-014
Cn3an12a1 TDn3a1 TDn12a1 2e-014
Cn3an12a2 TDn3a3 TDn12a3 1e-014
Cn3an12a3 TDn3a5 TDn12a5 1e-014
Cn3an12a4 TDn3a7 TDn12a7 1e-014
Cn3an12a5 TDn3a9 TDn12a9 1e-014
Cn3an12a6 TDn3a11 TDn12a11 1e-014
Cn3an12a7 TDn3a13 TDn12a13 1e-014
Cn3an12a8 TDn3a15 TDn12a15 1e-014
Cn3an12a9 TDn3a17 TDn12a17 1e-014
Cn3an12a10 TDn3a19 TDn12a19 1e-014
Cn3an12a11 TDn3a21 TDn12a21 1e-014
Cn3an12a12 TDn3a23 TDn12a23 1e-014
Cn3an12a13 TDn3a25 TDn12a25 1e-014
Cn3an12a14 TDn3a27 TDn12a27 1e-014
Cn3an12a15 TDn3a29 TDn12a29 1e-014
Cn3an12a16 TDn3a31 TDn12a31 1e-014
Cn3an12a17 TDn3a33 TDn12a33 2e-014
Cn3anva1 TDn3a1 TDnva1 2e-014
Cn3anva2 TDn3a3 TDnva3 2e-014
Cn3anva3 TDn3a5 TDnva5 2e-014
Cn3anva4 TDn3a7 TDnva7 2e-014
Cn3anva5 TDn3a9 TDnva9 2e-014
Cn3anva6 TDn3a11 TDnva11 2e-014
Cn3anva7 TDn3a13 TDnva13 2e-014
Cn3anva8 TDn3a15 TDnva15 2e-014
Cn3anva9 TDn3a17 TDnva17 2e-014
Cn3anva10 TDn3a19 TDnva19 2e-014
Cn3anva11 TDn3a21 TDnva21 2e-014
Cn3anva12 TDn3a23 TDnva23 2e-014
Cn3anva13 TDn3a25 TDnva25 2e-014
Cn3anva14 TDn3a27 TDnva27 2e-014
Cn3anva15 TDn3a29 TDnva29 2e-014
Cn3anva16 TDn3a31 TDnva31 2e-014
Cn3anva17 TDn3a33 TDnva33 2e-014
Cn4an5a1 TDn4a1 TDn5a1 1.573240e-014
Cn4an5a2 TDn4a3 TDn5a3 3e-014
Cn4an5a3 TDn4a5 TDn5a5 3e-014
Cn4an5a4 TDn4a7 TDn5a7 3e-014
Cn4an5a5 TDn4a9 TDn5a9 3e-014
Cn4an5a6 TDn4a11 TDn5a11 3e-014
Cn4an5a7 TDn4a13 TDn5a13 3e-014
Cn4an5a8 TDn4a15 TDn5a15 3e-014
Cn4an5a9 TDn4a17 TDn5a17 3e-014
Cn4an5a10 TDn4a19 TDn5a19 3e-014
Cn4an5a11 TDn4a21 TDn5a21 3e-014
Cn4an5a12 TDn4a23 TDn5a23 3e-014
Cn4an5a13 TDn4a25 TDn5a25 3e-014
Cn4an5a14 TDn4a27 TDn5a27 3e-014
Cn4an5a15 TDn4a29 TDn5a29 3e-014
Cn4an5a16 TDn4a31 TDn5a31 3e-014
Cn4an5a17 TDn4a33 TDn5a33 1.573240e-014
Cn4an6a1 TDn4a1 TDn6a1 5.586810e-015
Cn4an6a2 TDn4a3 TDn6a3 1e-014
Cn4an6a3 TDn4a5 TDn6a5 1e-014
Cn4an6a4 TDn4a7 TDn6a7 1e-014
Cn4an6a5 TDn4a9 TDn6a9 1e-014
Cn4an6a6 TDn4a11 TDn6a11 1e-014
Cn4an6a7 TDn4a13 TDn6a13 1e-014
Cn4an6a8 TDn4a15 TDn6a15 1e-014
Cn4an6a9 TDn4a17 TDn6a17 1e-014
Cn4an6a10 TDn4a19 TDn6a19 1e-014
Cn4an6a11 TDn4a21 TDn6a21 1e-014
Cn4an6a12 TDn4a23 TDn6a23 1e-014
Cn4an6a13 TDn4a25 TDn6a25 1e-014
Cn4an6a14 TDn4a27 TDn6a27 1e-014
Cn4an6a15 TDn4a29 TDn6a29 1e-014
Cn4an6a16 TDn4a31 TDn6a31 1e-014
Cn4an6a17 TDn4a33 TDn6a33 5.586810e-015
Cn4an7a1 TDn4a1 TDn7a1 5.148610e-015
Cn4an7a2 TDn4a3 TDn7a3 1e-014
Cn4an7a3 TDn4a5 TDn7a5 1e-014
Cn4an7a4 TDn4a7 TDn7a7 1e-014
Cn4an7a5 TDn4a9 TDn7a9 1e-014
Cn4an7a6 TDn4a11 TDn7a11 1e-014
Cn4an7a7 TDn4a13 TDn7a13 1e-014
Cn4an7a8 TDn4a15 TDn7a15 1e-014
Cn4an7a9 TDn4a17 TDn7a17 1e-014
Cn4an7a10 TDn4a19 TDn7a19 1e-014
Cn4an7a11 TDn4a21 TDn7a21 1e-014
Cn4an7a12 TDn4a23 TDn7a23 1e-014
Cn4an7a13 TDn4a25 TDn7a25 1e-014
Cn4an7a14 TDn4a27 TDn7a27 1e-014
Cn4an7a15 TDn4a29 TDn7a29 1e-014
Cn4an7a16 TDn4a31 TDn7a31 1e-014
Cn4an7a17 TDn4a33 TDn7a33 5.148610e-015
Cn4an8a1 TDn4a1 TDn8a1 5.060570e-015
Cn4an8a2 TDn4a3 TDn8a3 1e-014
Cn4an8a3 TDn4a5 TDn8a5 1e-014
Cn4an8a4 TDn4a7 TDn8a7 1e-014
Cn4an8a5 TDn4a9 TDn8a9 1e-014
Cn4an8a6 TDn4a11 TDn8a11 1e-014
Cn4an8a7 TDn4a13 TDn8a13 1e-014
Cn4an8a8 TDn4a15 TDn8a15 1e-014
Cn4an8a9 TDn4a17 TDn8a17 1e-014
Cn4an8a10 TDn4a19 TDn8a19 1e-014
Cn4an8a11 TDn4a21 TDn8a21 1e-014
Cn4an8a12 TDn4a23 TDn8a23 1e-014
Cn4an8a13 TDn4a25 TDn8a25 1e-014
Cn4an8a14 TDn4a27 TDn8a27 1e-014
Cn4an8a15 TDn4a29 TDn8a29 1e-014
Cn4an8a16 TDn4a31 TDn8a31 1e-014
Cn4an8a17 TDn4a33 TDn8a33 5.060570e-015
Cn4an9a1 TDn4a1 TDn9a1 5.736010e-015
Cn4an9a2 TDn4a3 TDn9a3 1e-014
Cn4an9a3 TDn4a5 TDn9a5 1e-014
Cn4an9a4 TDn4a7 TDn9a7 1e-014
Cn4an9a5 TDn4a9 TDn9a9 1e-014
Cn4an9a6 TDn4a11 TDn9a11 1e-014
Cn4an9a7 TDn4a13 TDn9a13 1e-014
Cn4an9a8 TDn4a15 TDn9a15 1e-014
Cn4an9a9 TDn4a17 TDn9a17 1e-014
Cn4an9a10 TDn4a19 TDn9a19 1e-014
Cn4an9a11 TDn4a21 TDn9a21 1e-014
Cn4an9a12 TDn4a23 TDn9a23 1e-014
Cn4an9a13 TDn4a25 TDn9a25 1e-014
Cn4an9a14 TDn4a27 TDn9a27 1e-014
Cn4an9a15 TDn4a29 TDn9a29 1e-014
Cn4an9a16 TDn4a31 TDn9a31 1e-014
Cn4an9a17 TDn4a33 TDn9a33 5.736010e-015
Cn4an10a1 TDn4a1 TDn10a1 2e-014
Cn4an10a2 TDn4a3 TDn10a3 1e-014
Cn4an10a3 TDn4a5 TDn10a5 1e-014
Cn4an10a4 TDn4a7 TDn10a7 1e-014
Cn4an10a5 TDn4a9 TDn10a9 1e-014
Cn4an10a6 TDn4a11 TDn10a11 1e-014
Cn4an10a7 TDn4a13 TDn10a13 1e-014
Cn4an10a8 TDn4a15 TDn10a15 1e-014
Cn4an10a9 TDn4a17 TDn10a17 1e-014
Cn4an10a10 TDn4a19 TDn10a19 1e-014
Cn4an10a11 TDn4a21 TDn10a21 1e-014
Cn4an10a12 TDn4a23 TDn10a23 1e-014
Cn4an10a13 TDn4a25 TDn10a25 1e-014
Cn4an10a14 TDn4a27 TDn10a27 1e-014
Cn4an10a15 TDn4a29 TDn10a29 1e-014
Cn4an10a16 TDn4a31 TDn10a31 1e-014
Cn4an10a17 TDn4a33 TDn10a33 2e-014
Cn4an11a1 TDn4a1 TDn11a1 2e-014
Cn4an11a2 TDn4a3 TDn11a3 1e-014
Cn4an11a3 TDn4a5 TDn11a5 1e-014
Cn4an11a4 TDn4a7 TDn11a7 1e-014
Cn4an11a5 TDn4a9 TDn11a9 1e-014
Cn4an11a6 TDn4a11 TDn11a11 1e-014
Cn4an11a7 TDn4a13 TDn11a13 1e-014
Cn4an11a8 TDn4a15 TDn11a15 1e-014
Cn4an11a9 TDn4a17 TDn11a17 1e-014
Cn4an11a10 TDn4a19 TDn11a19 1e-014
Cn4an11a11 TDn4a21 TDn11a21 1e-014
Cn4an11a12 TDn4a23 TDn11a23 1e-014
Cn4an11a13 TDn4a25 TDn11a25 1e-014
Cn4an11a14 TDn4a27 TDn11a27 1e-014
Cn4an11a15 TDn4a29 TDn11a29 1e-014
Cn4an11a16 TDn4a31 TDn11a31 1e-014
Cn4an11a17 TDn4a33 TDn11a33 2e-014
Cn4an12a1 TDn4a1 TDn12a1 2e-014
Cn4an12a2 TDn4a3 TDn12a3 1e-014
Cn4an12a3 TDn4a5 TDn12a5 1e-014
Cn4an12a4 TDn4a7 TDn12a7 1e-014
Cn4an12a5 TDn4a9 TDn12a9 1e-014
Cn4an12a6 TDn4a11 TDn12a11 1e-014
Cn4an12a7 TDn4a13 TDn12a13 1e-014
Cn4an12a8 TDn4a15 TDn12a15 1e-014
Cn4an12a9 TDn4a17 TDn12a17 1e-014
Cn4an12a10 TDn4a19 TDn12a19 1e-014
Cn4an12a11 TDn4a21 TDn12a21 1e-014
Cn4an12a12 TDn4a23 TDn12a23 1e-014
Cn4an12a13 TDn4a25 TDn12a25 1e-014
Cn4an12a14 TDn4a27 TDn12a27 1e-014
Cn4an12a15 TDn4a29 TDn12a29 1e-014
Cn4an12a16 TDn4a31 TDn12a31 1e-014
Cn4an12a17 TDn4a33 TDn12a33 2e-014
Cn4anva1 TDn4a1 TDnva1 2e-014
Cn4anva2 TDn4a3 TDnva3 2e-014
Cn4anva3 TDn4a5 TDnva5 2e-014
Cn4anva4 TDn4a7 TDnva7 2e-014
Cn4anva5 TDn4a9 TDnva9 2e-014
Cn4anva6 TDn4a11 TDnva11 2e-014
Cn4anva7 TDn4a13 TDnva13 2e-014
Cn4anva8 TDn4a15 TDnva15 2e-014
Cn4anva9 TDn4a17 TDnva17 2e-014
Cn4anva10 TDn4a19 TDnva19 2e-014
Cn4anva11 TDn4a21 TDnva21 2e-014
Cn4anva12 TDn4a23 TDnva23 2e-014
Cn4anva13 TDn4a25 TDnva25 2e-014
Cn4anva14 TDn4a27 TDnva27 2e-014
Cn4anva15 TDn4a29 TDnva29 2e-014
Cn4anva16 TDn4a31 TDnva31 2e-014
Cn4anva17 TDn4a33 TDnva33 2e-014
Cn5an6a1 TDn5a1 TDn6a1 1.575710e-014
Cn5an6a2 TDn5a3 TDn6a3 3e-014
Cn5an6a3 TDn5a5 TDn6a5 3e-014
Cn5an6a4 TDn5a7 TDn6a7 3e-014
Cn5an6a5 TDn5a9 TDn6a9 3e-014
Cn5an6a6 TDn5a11 TDn6a11 3e-014
Cn5an6a7 TDn5a13 TDn6a13 3e-014
Cn5an6a8 TDn5a15 TDn6a15 3e-014
Cn5an6a9 TDn5a17 TDn6a17 3e-014
Cn5an6a10 TDn5a19 TDn6a19 3e-014
Cn5an6a11 TDn5a21 TDn6a21 3e-014
Cn5an6a12 TDn5a23 TDn6a23 3e-014
Cn5an6a13 TDn5a25 TDn6a25 3e-014
Cn5an6a14 TDn5a27 TDn6a27 3e-014
Cn5an6a15 TDn5a29 TDn6a29 3e-014
Cn5an6a16 TDn5a31 TDn6a31 3e-014
Cn5an6a17 TDn5a33 TDn6a33 1.575710e-014
Cn5an7a1 TDn5a1 TDn7a1 5.608560e-015
Cn5an7a2 TDn5a3 TDn7a3 1e-014
Cn5an7a3 TDn5a5 TDn7a5 1e-014
Cn5an7a4 TDn5a7 TDn7a7 1e-014
Cn5an7a5 TDn5a9 TDn7a9 1e-014
Cn5an7a6 TDn5a11 TDn7a11 1e-014
Cn5an7a7 TDn5a13 TDn7a13 1e-014
Cn5an7a8 TDn5a15 TDn7a15 1e-014
Cn5an7a9 TDn5a17 TDn7a17 1e-014
Cn5an7a10 TDn5a19 TDn7a19 1e-014
Cn5an7a11 TDn5a21 TDn7a21 1e-014
Cn5an7a12 TDn5a23 TDn7a23 1e-014
Cn5an7a13 TDn5a25 TDn7a25 1e-014
Cn5an7a14 TDn5a27 TDn7a27 1e-014
Cn5an7a15 TDn5a29 TDn7a29 1e-014
Cn5an7a17 TDn5a33 TDn7a33 5.608560e-015
Cn5an8a1 TDn5a1 TDn8a1 5.204690e-015
Cn5an8a2 TDn5a3 TDn8a3 1e-014
Cn5an8a3 TDn5a5 TDn8a5 1e-014
Cn5an8a4 TDn5a7 TDn8a7 1e-014
Cn5an8a5 TDn5a9 TDn8a9 1e-014
Cn5an8a6 TDn5a11 TDn8a11 1e-014
Cn5an8a7 TDn5a13 TDn8a13 1e-014
Cn5an8a8 TDn5a15 TDn8a15 1e-014
Cn5an8a9 TDn5a17 TDn8a17 1e-014
Cn5an8a10 TDn5a19 TDn8a19 1e-014
Cn5an8a11 TDn5a21 TDn8a21 1e-014
Cn5an8a12 TDn5a23 TDn8a23 1e-014
Cn5an8a13 TDn5a25 TDn8a25 1e-014
Cn5an8a14 TDn5a27 TDn8a27 1e-014
Cn5an8a15 TDn5a29 TDn8a29 1e-014
Cn5an8a16 TDn5a31 TDn8a31 1e-014
Cn5an8a17 TDn5a33 TDn8a33 5.204690e-015
Cn5an9a1 TDn5a1 TDn9a1 5.818520e-015
Cn5an9a2 TDn5a3 TDn9a3 1e-014
Cn5an9a3 TDn5a5 TDn9a5 1e-014
Cn5an9a4 TDn5a7 TDn9a7 1e-014
Cn5an9a5 TDn5a9 TDn9a9 1e-014
Cn5an9a6 TDn5a11 TDn9a11 1e-014
Cn5an9a7 TDn5a13 TDn9a13 1e-014
Cn5an9a8 TDn5a15 TDn9a15 1e-014
Cn5an9a9 TDn5a17 TDn9a17 1e-014
Cn5an9a10 TDn5a19 TDn9a19 1e-014
Cn5an9a11 TDn5a21 TDn9a21 1e-014
Cn5an9a12 TDn5a23 TDn9a23 1e-014
Cn5an9a13 TDn5a25 TDn9a25 1e-014
Cn5an9a14 TDn5a27 TDn9a27 1e-014
Cn5an9a15 TDn5a29 TDn9a29 1e-014
Cn5an9a16 TDn5a31 TDn9a31 1e-014
Cn5an9a17 TDn5a33 TDn9a33 5.818520e-015
Cn5an10a1 TDn5a1 TDn10a1 2e-014
Cn5an10a2 TDn5a3 TDn10a3 1e-014
Cn5an10a3 TDn5a5 TDn10a5 1e-014
Cn5an10a4 TDn5a7 TDn10a7 1e-014
Cn5an10a5 TDn5a9 TDn10a9 1e-014
Cn5an10a6 TDn5a11 TDn10a11 1e-014
Cn5an10a7 TDn5a13 TDn10a13 1e-014
Cn5an10a8 TDn5a15 TDn10a15 1e-014
Cn5an10a9 TDn5a17 TDn10a17 1e-014
Cn5an10a10 TDn5a19 TDn10a19 1e-014
Cn5an10a11 TDn5a21 TDn10a21 1e-014
Cn5an10a12 TDn5a23 TDn10a23 1e-014
Cn5an10a13 TDn5a25 TDn10a25 1e-014
Cn5an10a14 TDn5a27 TDn10a27 1e-014
Cn5an10a15 TDn5a29 TDn10a29 1e-014
Cn5an10a16 TDn5a31 TDn10a31 1e-014
Cn5an10a17 TDn5a33 TDn10a33 2e-014
Cn5an11a1 TDn5a1 TDn11a1 2e-014
Cn5an11a2 TDn5a3 TDn11a3 1e-014
Cn5an11a3 TDn5a5 TDn11a5 1e-014
Cn5an11a4 TDn5a7 TDn11a7 1e-014
Cn5an11a5 TDn5a9 TDn11a9 1e-014
Cn5an11a6 TDn5a11 TDn11a11 1e-014
Cn5an11a7 TDn5a13 TDn11a13 1e-014
Cn5an11a8 TDn5a15 TDn11a15 1e-014
Cn5an11a9 TDn5a17 TDn11a17 1e-014
Cn5an11a10 TDn5a19 TDn11a19 1e-014
Cn5an11a11 TDn5a21 TDn11a21 1e-014
Cn5an11a12 TDn5a23 TDn11a23 1e-014
Cn5an11a13 TDn5a25 TDn11a25 1e-014
Cn5an11a14 TDn5a27 TDn11a27 1e-014
Cn5an11a15 TDn5a29 TDn11a29 1e-014
Cn5an11a16 TDn5a31 TDn11a31 1e-014
Cn5an11a17 TDn5a33 TDn11a33 2e-014
Cn5an12a1 TDn5a1 TDn12a1 2e-014
Cn5an12a2 TDn5a3 TDn12a3 1e-014
Cn5an12a3 TDn5a5 TDn12a5 1e-014
Cn5an12a4 TDn5a7 TDn12a7 1e-014
Cn5an12a5 TDn5a9 TDn12a9 1e-014
Cn5an12a6 TDn5a11 TDn12a11 1e-014
Cn5an12a7 TDn5a13 TDn12a13 1e-014
Cn5an12a8 TDn5a15 TDn12a15 1e-014
Cn5an12a9 TDn5a17 TDn12a17 1e-014
Cn5an12a10 TDn5a19 TDn12a19 1e-014
Cn5an12a11 TDn5a21 TDn12a21 1e-014
Cn5an12a12 TDn5a23 TDn12a23 1e-014
Cn5an12a13 TDn5a25 TDn12a25 1e-014
Cn5an12a14 TDn5a27 TDn12a27 1e-014
Cn5an12a15 TDn5a29 TDn12a29 1e-014
Cn5an12a16 TDn5a31 TDn12a31 1e-014
Cn5an12a17 TDn5a33 TDn12a33 2e-014
Cn5anva1 TDn5a1 TDnva1 2e-014
Cn5anva2 TDn5a3 TDnva3 2e-014
Cn5anva3 TDn5a5 TDnva5 2e-014
Cn5anva4 TDn5a7 TDnva7 2e-014
Cn5anva5 TDn5a9 TDnva9 2e-014
Cn5anva6 TDn5a11 TDnva11 2e-014
Cn5anva7 TDn5a13 TDnva13 2e-014
Cn5anva8 TDn5a15 TDnva15 2e-014
Cn5anva9 TDn5a17 TDnva17 2e-014
Cn5anva10 TDn5a19 TDnva19 2e-014
Cn5anva11 TDn5a21 TDnva21 2e-014
Cn5anva12 TDn5a23 TDnva23 2e-014
Cn5anva13 TDn5a25 TDnva25 2e-014
Cn5anva14 TDn5a27 TDnva27 2e-014
Cn5anva15 TDn5a29 TDnva29 2e-014
Cn5anva16 TDn5a31 TDnva31 2e-014
Cn5anva17 TDn5a33 TDnva33 2e-014
Cn6an7a1 TDn6a1 TDn7a1 1.578870e-014
Cn6an7a2 TDn6a3 TDn7a3 3e-014
Cn6an7a3 TDn6a5 TDn7a5 3e-014
Cn6an7a4 TDn6a7 TDn7a7 3e-014
Cn6an7a5 TDn6a9 TDn7a9 3e-014
Cn6an7a6 TDn6a11 TDn7a11 3e-014
Cn6an7a7 TDn6a13 TDn7a13 3e-014
Cn6an7a8 TDn6a15 TDn7a15 3e-014
Cn6an7a9 TDn6a17 TDn7a17 3e-014
Cn6an7a10 TDn6a19 TDn7a19 3e-014
Cn6an7a11 TDn6a21 TDn7a21 3e-014
Cn6an7a12 TDn6a23 TDn7a23 3e-014
Cn6an7a13 TDn6a25 TDn7a25 3e-014
Cn6an7a14 TDn6a27 TDn7a27 3e-014
Cn6an7a15 TDn6a29 TDn7a29 3e-014
Cn6an7a16 TDn6a31 TDn7a31 3e-014
Cn6an7a17 TDn6a33 TDn7a33 1.578870e-014
Cn6an8a1 TDn6a1 TDn8a1 5.673080e-015
Cn6an8a2 TDn6a3 TDn8a3 1e-014
Cn6an8a3 TDn6a5 TDn8a5 1e-014
Cn6an8a4 TDn6a7 TDn8a7 1e-014
Cn6an8a5 TDn6a9 TDn8a9 1e-014
Cn6an8a6 TDn6a11 TDn8a11 1e-014
Cn6an8a7 TDn6a13 TDn8a13 1e-014
Cn6an8a8 TDn6a15 TDn8a15 1e-014
Cn6an8a9 TDn6a17 TDn8a17 1e-014
Cn6an8a10 TDn6a19 TDn8a19 1e-014
Cn6an8a11 TDn6a21 TDn8a21 1e-014
Cn6an8a12 TDn6a23 TDn8a23 1e-014
Cn6an8a13 TDn6a25 TDn8a25 1e-014
Cn6an8a14 TDn6a27 TDn8a27 1e-014
Cn6an8a15 TDn6a29 TDn8a29 1e-014
Cn6an8a16 TDn6a31 TDn8a31 1e-014
Cn6an8a17 TDn6a33 TDn8a33 5.673080e-015
Cn6an9a1 TDn6a1 TDn9a1 6.001130e-015
Cn6an9a2 TDn6a3 TDn9a3 1e-014
Cn6an9a3 TDn6a5 TDn9a5 1e-014
Cn6an9a4 TDn6a7 TDn9a7 1e-014
Cn6an9a5 TDn6a9 TDn9a9 1e-014
Cn6an9a6 TDn6a11 TDn9a11 1e-014
Cn6an9a7 TDn6a13 TDn9a13 1e-014
Cn6an9a8 TDn6a15 TDn9a15 1e-014
Cn6an9a9 TDn6a17 TDn9a17 1e-014
Cn6an9a10 TDn6a19 TDn9a19 1e-014
Cn6an9a11 TDn6a21 TDn9a21 1e-014
Cn6an9a12 TDn6a23 TDn9a23 1e-014
Cn6an9a13 TDn6a25 TDn9a25 1e-014
Cn6an9a14 TDn6a27 TDn9a27 1e-014
Cn6an9a15 TDn6a29 TDn9a29 1e-014
Cn6an9a16 TDn6a31 TDn9a31 1e-014
Cn6an9a17 TDn6a33 TDn9a33 6.001130e-015
Cn6an10a1 TDn6a1 TDn10a1 2e-014
Cn6an10a2 TDn6a3 TDn10a3 1e-014
Cn6an10a3 TDn6a5 TDn10a5 1e-014
Cn6an10a4 TDn6a7 TDn10a7 1e-014
Cn6an10a5 TDn6a9 TDn10a9 1e-014
Cn6an10a6 TDn6a11 TDn10a11 1e-014
Cn6an10a7 TDn6a13 TDn10a13 1e-014
Cn6an10a8 TDn6a15 TDn10a15 1e-014
Cn6an10a9 TDn6a17 TDn10a17 1e-014
Cn6an10a10 TDn6a19 TDn10a19 1e-014
Cn6an10a11 TDn6a21 TDn10a21 1e-014
Cn6an10a12 TDn6a23 TDn10a23 1e-014
Cn6an10a13 TDn6a25 TDn10a25 1e-014
Cn6an10a14 TDn6a27 TDn10a27 1e-014
Cn6an10a15 TDn6a29 TDn10a29 1e-014
Cn6an10a16 TDn6a31 TDn10a31 1e-014
Cn6an10a17 TDn6a33 TDn10a33 2e-014
Cn6an11a1 TDn6a1 TDn11a1 2e-014
Cn6an11a2 TDn6a3 TDn11a3 1e-014
Cn6an11a3 TDn6a5 TDn11a5 1e-014
Cn6an11a4 TDn6a7 TDn11a7 1e-014
Cn6an11a5 TDn6a9 TDn11a9 1e-014
Cn6an11a6 TDn6a11 TDn11a11 1e-014
Cn6an11a7 TDn6a13 TDn11a13 1e-014
Cn6an11a8 TDn6a15 TDn11a15 1e-014
Cn6an11a9 TDn6a17 TDn11a17 1e-014
Cn6an11a10 TDn6a19 TDn11a19 1e-014
Cn6an11a11 TDn6a21 TDn11a21 1e-014
Cn6an11a12 TDn6a23 TDn11a23 1e-014
Cn6an11a13 TDn6a25 TDn11a25 1e-014
Cn6an11a14 TDn6a27 TDn11a27 1e-014
Cn6an11a15 TDn6a29 TDn11a29 1e-014
Cn6an11a16 TDn6a31 TDn11a31 1e-014
Cn6an11a17 TDn6a33 TDn11a33 2e-014
Cn6an12a1 TDn6a1 TDn12a1 2e-014
Cn6an12a2 TDn6a3 TDn12a3 1e-014
Cn6an12a3 TDn6a5 TDn12a5 1e-014
Cn6an12a4 TDn6a7 TDn12a7 1e-014
Cn6an12a5 TDn6a9 TDn12a9 1e-014
Cn6an12a6 TDn6a11 TDn12a11 1e-014
Cn6an12a7 TDn6a13 TDn12a13 1e-014
Cn6an12a8 TDn6a15 TDn12a15 1e-014
Cn6an12a9 TDn6a17 TDn12a17 1e-014
Cn6an12a10 TDn6a19 TDn12a19 1e-014
Cn6an12a11 TDn6a21 TDn12a21 1e-014
Cn6an12a12 TDn6a23 TDn12a23 1e-014
Cn6an12a13 TDn6a25 TDn12a25 1e-014
Cn6an12a14 TDn6a27 TDn12a27 1e-014
Cn6an12a15 TDn6a29 TDn12a29 1e-014
Cn6an12a16 TDn6a31 TDn12a31 1e-014
Cn6an12a17 TDn6a33 TDn12a33 2e-014
Cn6anva1 TDn6a1 TDnva1 2e-014
Cn6anva2 TDn6a3 TDnva3 2e-014
Cn6anva3 TDn6a5 TDnva5 2e-014
Cn6anva4 TDn6a7 TDnva7 2e-014
Cn6anva5 TDn6a9 TDnva9 2e-014
Cn6anva6 TDn6a11 TDnva11 2e-014
Cn6anva7 TDn6a13 TDnva13 2e-014
Cn6anva8 TDn6a15 TDnva15 2e-014
Cn6anva9 TDn6a17 TDnva17 2e-014
Cn6anva10 TDn6a19 TDnva19 2e-014
Cn6anva11 TDn6a21 TDnva21 2e-014
Cn6anva12 TDn6a23 TDnva23 2e-014
Cn6anva13 TDn6a25 TDnva25 2e-014
Cn6anva14 TDn6a27 TDnva27 2e-014
Cn6anva15 TDn6a29 TDnva29 2e-014
Cn6anva16 TDn6a31 TDnva31 2e-014
Cn6anva17 TDn6a33 TDnva33 2e-014
Cn7an8a1 TDn7a1 TDn8a1 1.587490e-014
Cn7an8a2 TDn7a3 TDn8a3 3e-014
Cn7an8a3 TDn7a5 TDn8a5 3e-014
Cn7an8a4 TDn7a7 TDn8a7 3e-014
Cn7an8a5 TDn7a9 TDn8a9 3e-014
Cn7an8a6 TDn7a11 TDn8a11 3e-014
Cn7an8a7 TDn7a13 TDn8a13 3e-014
Cn7an8a8 TDn7a15 TDn8a15 3e-014
Cn7an8a9 TDn7a17 TDn8a17 3e-014
Cn7an8a10 TDn7a19 TDn8a19 3e-014
Cn7an8a11 TDn7a21 TDn8a21 3e-014
Cn7an8a12 TDn7a23 TDn8a23 3e-014
Cn7an8a13 TDn7a25 TDn8a25 3e-014
Cn7an8a14 TDn7a27 TDn8a27 3e-014
Cn7an8a15 TDn7a29 TDn8a29 3e-014
Cn7an8a16 TDn7a31 TDn8a31 3e-014
Cn7an8a17 TDn7a33 TDn8a33 1.587490e-014
Cn7an9a1 TDn7a1 TDn9a1 6.511580e-015
Cn7an9a2 TDn7a3 TDn9a3 1e-014
Cn7an9a3 TDn7a5 TDn9a5 1e-014
Cn7an9a4 TDn7a7 TDn9a7 1e-014
Cn7an9a5 TDn7a9 TDn9a9 1e-014
Cn7an9a6 TDn7a11 TDn9a11 1e-014
Cn7an9a7 TDn7a13 TDn9a13 1e-014
Cn7an9a8 TDn7a15 TDn9a15 1e-014
Cn7an9a9 TDn7a17 TDn9a17 1e-014
Cn7an9a10 TDn7a19 TDn9a19 1e-014
Cn7an9a11 TDn7a21 TDn9a21 1e-014
Cn7an9a12 TDn7a23 TDn9a23 1e-014
Cn7an9a13 TDn7a25 TDn9a25 1e-014
Cn7an9a14 TDn7a27 TDn9a27 1e-014
Cn7an9a15 TDn7a29 TDn9a29 1e-014
Cn7an9a16 TDn7a31 TDn9a31 1e-014
Cn7an9a17 TDn7a33 TDn9a33 6.511580e-015
Cn7an10a1 TDn7a1 TDn10a1 2e-014
Cn7an10a2 TDn7a3 TDn10a3 1e-014
Cn7an10a3 TDn7a5 TDn10a5 1e-014
Cn7an10a4 TDn7a7 TDn10a7 1e-014
Cn7an10a5 TDn7a9 TDn10a9 1e-014
Cn7an10a6 TDn7a11 TDn10a11 1e-014
Cn7an10a7 TDn7a13 TDn10a13 1e-014
Cn7an10a8 TDn7a15 TDn10a15 1e-014
Cn7an10a9 TDn7a17 TDn10a17 1e-014
Cn7an10a10 TDn7a19 TDn10a19 1e-014
Cn7an10a11 TDn7a21 TDn10a21 1e-014
Cn7an10a12 TDn7a23 TDn10a23 1e-014
Cn7an10a13 TDn7a25 TDn10a25 1e-014
Cn7an10a14 TDn7a27 TDn10a27 1e-014
Cn7an10a15 TDn7a29 TDn10a29 1e-014
Cn7an10a16 TDn7a31 TDn10a31 1e-014
Cn7an10a17 TDn7a33 TDn10a33 2e-014
Cn7an11a1 TDn7a1 TDn11a1 2e-014
Cn7an11a2 TDn7a3 TDn11a3 1e-014
Cn7an11a3 TDn7a5 TDn11a5 1e-014
Cn7an11a4 TDn7a7 TDn11a7 1e-014
Cn7an11a5 TDn7a9 TDn11a9 1e-014
Cn7an11a6 TDn7a11 TDn11a11 1e-014
Cn7an11a7 TDn7a13 TDn11a13 1e-014
Cn7an11a8 TDn7a15 TDn11a15 1e-014
Cn7an11a9 TDn7a17 TDn11a17 1e-014
Cn7an11a10 TDn7a19 TDn11a19 1e-014
Cn7an11a11 TDn7a21 TDn11a21 1e-014
Cn7an11a12 TDn7a23 TDn11a23 1e-014
Cn7an11a13 TDn7a25 TDn11a25 1e-014
Cn7an11a14 TDn7a27 TDn11a27 1e-014
Cn7an11a15 TDn7a29 TDn11a29 1e-014
Cn7an11a16 TDn7a31 TDn11a31 1e-014
Cn7an11a17 TDn7a33 TDn11a33 2e-014
Cn7an12a1 TDn7a1 TDn12a1 2e-014
Cn7an12a2 TDn7a3 TDn12a3 1e-014
Cn7an12a3 TDn7a5 TDn12a5 1e-014
Cn7an12a4 TDn7a7 TDn12a7 1e-014
Cn7an12a5 TDn7a9 TDn12a9 1e-014
Cn7an12a6 TDn7a11 TDn12a11 1e-014
Cn7an12a7 TDn7a13 TDn12a13 1e-014
Cn7an12a8 TDn7a15 TDn12a15 1e-014
Cn7an12a9 TDn7a17 TDn12a17 1e-014
Cn7an12a10 TDn7a19 TDn12a19 1e-014
Cn7an12a11 TDn7a21 TDn12a21 1e-014
Cn7an12a12 TDn7a23 TDn12a23 1e-014
Cn7an12a13 TDn7a25 TDn12a25 1e-014
Cn7an12a14 TDn7a27 TDn12a27 1e-014
Cn7an12a15 TDn7a29 TDn12a29 1e-014
Cn7an12a16 TDn7a31 TDn12a31 1e-014
Cn7an12a17 TDn7a33 TDn12a33 2e-014
Cn7anva1 TDn7a1 TDnva1 2e-014
Cn7anva2 TDn7a3 TDnva3 2e-014
Cn7anva3 TDn7a5 TDnva5 2e-014
Cn7anva4 TDn7a7 TDnva7 2e-014
Cn7anva5 TDn7a9 TDnva9 2e-014
Cn7anva6 TDn7a11 TDnva11 2e-014
Cn7anva7 TDn7a13 TDnva13 2e-014
Cn7anva8 TDn7a15 TDnva15 2e-014
Cn7anva9 TDn7a17 TDnva17 2e-014
Cn7anva10 TDn7a19 TDnva19 2e-014
Cn7anva11 TDn7a21 TDnva21 2e-014
Cn7anva12 TDn7a23 TDnva23 2e-014
Cn7anva13 TDn7a25 TDnva25 2e-014
Cn7anva14 TDn7a27 TDnva27 2e-014
Cn7anva15 TDn7a29 TDnva29 2e-014
Cn7anva16 TDn7a31 TDnva31 2e-014
Cn7anva17 TDn7a33 TDnva33 2e-014
Cn8an9a1 TDn8a1 TDn9a1 2e-014
Cn8an9a2 TDn8a3 TDn9a3 3e-014
Cn8an9a3 TDn8a5 TDn9a5 3e-014
Cn8an9a4 TDn8a7 TDn9a7 3e-014
Cn8an9a5 TDn8a9 TDn9a9 3e-014
Cn8an9a6 TDn8a11 TDn9a11 3e-014
Cn8an9a7 TDn8a13 TDn9a13 3e-014
Cn8an9a8 TDn8a15 TDn9a15 3e-014
Cn8an9a9 TDn8a17 TDn9a17 3e-014
Cn8an9a10 TDn8a19 TDn9a19 3e-014
Cn8an9a11 TDn8a21 TDn9a21 3e-014
Cn8an9a12 TDn8a23 TDn9a23 3e-014
Cn8an9a13 TDn8a25 TDn9a25 3e-014
Cn8an9a14 TDn8a27 TDn9a27 3e-014
Cn8an9a15 TDn8a29 TDn9a29 3e-014
Cn8an9a16 TDn8a31 TDn9a31 3e-014
Cn8an9a17 TDn8a33 TDn9a33 2e-014
Cn8an10a1 TDn8a1 TDn10a1 2e-014
Cn8an10a2 TDn8a3 TDn10a3 1e-014
Cn8an10a3 TDn8a5 TDn10a5 1e-014
Cn8an10a4 TDn8a7 TDn10a7 1e-014
Cn8an10a5 TDn8a9 TDn10a9 1e-014
Cn8an10a6 TDn8a11 TDn10a11 1e-014
Cn8an10a7 TDn8a13 TDn10a13 1e-014
Cn8an10a8 TDn8a15 TDn10a15 1e-014
Cn8an10a9 TDn8a17 TDn10a17 1e-014
Cn8an10a10 TDn8a19 TDn10a19 1e-014
Cn8an10a11 TDn8a21 TDn10a21 1e-014
Cn8an10a12 TDn8a23 TDn10a23 1e-014
Cn8an10a13 TDn8a25 TDn10a25 1e-014
Cn8an10a14 TDn8a27 TDn10a27 1e-014
Cn8an10a15 TDn8a29 TDn10a29 1e-014
Cn8an10a16 TDn8a31 TDn10a31 1e-014
Cn8an10a17 TDn8a33 TDn10a33 2e-014
Cn8an11a1 TDn8a1 TDn11a1 2e-014
Cn8an11a2 TDn8a3 TDn11a3 1e-014
Cn8an11a3 TDn8a5 TDn11a5 1e-014
Cn8an11a4 TDn8a7 TDn11a7 1e-014
Cn8an11a5 TDn8a9 TDn11a9 1e-014
Cn8an11a6 TDn8a11 TDn11a11 1e-014
Cn8an11a7 TDn8a13 TDn11a13 1e-014
Cn8an11a8 TDn8a15 TDn11a15 1e-014
Cn8an11a9 TDn8a17 TDn11a17 1e-014
Cn8an11a10 TDn8a19 TDn11a19 1e-014
Cn8an11a11 TDn8a21 TDn11a21 1e-014
Cn8an11a12 TDn8a23 TDn11a23 1e-014
Cn8an11a13 TDn8a25 TDn11a25 1e-014
Cn8an11a14 TDn8a27 TDn11a27 1e-014
Cn8an11a15 TDn8a29 TDn11a29 1e-014
Cn8an11a16 TDn8a31 TDn11a31 1e-014
Cn8an11a17 TDn8a33 TDn11a33 2e-014
Cn8an12a1 TDn8a1 TDn12a1 2e-014
Cn8an12a2 TDn8a3 TDn12a3 1e-014
Cn8an12a3 TDn8a5 TDn12a5 1e-014
Cn8an12a4 TDn8a7 TDn12a7 1e-014
Cn8an12a5 TDn8a9 TDn12a9 1e-014
Cn8an12a6 TDn8a11 TDn12a11 1e-014
Cn8an12a7 TDn8a13 TDn12a13 1e-014
Cn8an12a8 TDn8a15 TDn12a15 1e-014
Cn8an12a9 TDn8a17 TDn12a17 1e-014
Cn8an12a10 TDn8a19 TDn12a19 1e-014
Cn8an12a11 TDn8a21 TDn12a21 1e-014
Cn8an12a12 TDn8a23 TDn12a23 1e-014
Cn8an12a13 TDn8a25 TDn12a25 1e-014
Cn8an12a14 TDn8a27 TDn12a27 1e-014
Cn8an12a15 TDn8a29 TDn12a29 1e-014
Cn8an12a16 TDn8a31 TDn12a31 1e-014
Cn8an12a17 TDn8a33 TDn12a33 2e-014
Cn8anva1 TDn8a1 TDnva1 2e-014
Cn8anva2 TDn8a3 TDnva3 2e-014
Cn8anva3 TDn8a5 TDnva5 2e-014
Cn8anva4 TDn8a7 TDnva7 2e-014
Cn8anva5 TDn8a9 TDnva9 2e-014
Cn8anva6 TDn8a11 TDnva11 2e-014
Cn8anva7 TDn8a13 TDnva13 2e-014
Cn8anva8 TDn8a15 TDnva15 2e-014
Cn8anva9 TDn8a17 TDnva17 2e-014
Cn8anva10 TDn8a19 TDnva19 2e-014
Cn8anva11 TDn8a21 TDnva21 2e-014
Cn8anva12 TDn8a23 TDnva23 2e-014
Cn8anva13 TDn8a25 TDnva25 2e-014
Cn8anva14 TDn8a27 TDnva27 2e-014
Cn8anva15 TDn8a29 TDnva29 2e-014
Cn8anva16 TDn8a31 TDnva31 2e-014
Cn8anva17 TDn8a33 TDnva33 2e-014
Cn9an10a1 TDn9a1 TDn10a1 2e-014
Cn9an10a2 TDn9a3 TDn10a3 1e-014
Cn9an10a3 TDn9a5 TDn10a5 1e-014
Cn9an10a4 TDn9a7 TDn10a7 1e-014
Cn9an10a5 TDn9a9 TDn10a9 1e-014
Cn9an10a6 TDn9a11 TDn10a11 1e-014
Cn9an10a7 TDn9a13 TDn10a13 1e-014
Cn9an10a8 TDn9a15 TDn10a15 1e-014
Cn9an10a9 TDn9a17 TDn10a17 1e-014
Cn9an10a10 TDn9a19 TDn10a19 1e-014
Cn9an10a11 TDn9a21 TDn10a21 1e-014
Cn9an10a12 TDn9a23 TDn10a23 1e-014
Cn9an10a13 TDn9a25 TDn10a25 1e-014
Cn9an10a14 TDn9a27 TDn10a27 1e-014
Cn9an10a15 TDn9a29 TDn10a29 1e-014
Cn9an10a16 TDn9a31 TDn10a31 1e-014
Cn9an10a17 TDn9a33 TDn10a33 2e-014
Cn9an11a1 TDn9a1 TDn11a1 2e-014
Cn9an11a2 TDn9a3 TDn11a3 1e-014
Cn9an11a3 TDn9a5 TDn11a5 1e-014
Cn9an11a4 TDn9a7 TDn11a7 1e-014
Cn9an11a5 TDn9a9 TDn11a9 1e-014
Cn9an11a6 TDn9a11 TDn11a11 1e-014
Cn9an11a7 TDn9a13 TDn11a13 1e-014
Cn9an11a8 TDn9a15 TDn11a15 1e-014
Cn9an11a9 TDn9a17 TDn11a17 1e-014
Cn9an11a10 TDn9a19 TDn11a19 1e-014
Cn9an11a11 TDn9a21 TDn11a21 1e-014
Cn9an11a12 TDn9a23 TDn11a23 1e-014
Cn9an11a13 TDn9a25 TDn11a25 1e-014
Cn9an11a14 TDn9a27 TDn11a27 1e-014
Cn9an11a15 TDn9a29 TDn11a29 1e-014
Cn9an11a16 TDn9a31 TDn11a31 1e-014
Cn9an11a17 TDn9a33 TDn11a33 2e-014
Cn9an12a1 TDn9a1 TDn12a1 2e-014
Cn9an12a2 TDn9a3 TDn12a3 1e-014
Cn9an12a3 TDn9a5 TDn12a5 1e-014
Cn9an12a4 TDn9a7 TDn12a7 1e-014
Cn9an12a5 TDn9a9 TDn12a9 1e-014
Cn9an12a6 TDn9a11 TDn12a11 1e-014
Cn9an12a7 TDn9a13 TDn12a13 1e-014
Cn9an12a8 TDn9a15 TDn12a15 1e-014
Cn9an12a9 TDn9a17 TDn12a17 1e-014
Cn9an12a10 TDn9a19 TDn12a19 1e-014
Cn9an12a11 TDn9a21 TDn12a21 1e-014
Cn9an12a12 TDn9a23 TDn12a23 1e-014
Cn9an12a13 TDn9a25 TDn12a25 1e-014
Cn9an12a14 TDn9a27 TDn12a27 1e-014
Cn9an12a15 TDn9a29 TDn12a29 1e-014
Cn9an12a16 TDn9a31 TDn12a31 1e-014
Cn9an12a17 TDn9a33 TDn12a33 2e-014
Cn9anva1 TDn9a1 TDnva1 2e-014
Cn9anva2 TDn9a3 TDnva3 2e-014
Cn9anva3 TDn9a5 TDnva5 2e-014
Cn9anva4 TDn9a7 TDnva7 2e-014
Cn9anva5 TDn9a9 TDnva9 2e-014
Cn9anva6 TDn9a11 TDnva11 2e-014
Cn9anva7 TDn9a13 TDnva13 2e-014
Cn9anva8 TDn9a15 TDnva15 2e-014
Cn9anva9 TDn9a17 TDnva17 2e-014
Cn9anva10 TDn9a19 TDnva19 2e-014
Cn9anva11 TDn9a21 TDnva21 2e-014
Cn9anva12 TDn9a23 TDnva23 2e-014
Cn9anva13 TDn9a25 TDnva25 2e-014
Cn9anva14 TDn9a27 TDnva27 2e-014
Cn9anva15 TDn9a29 TDnva29 2e-014
Cn9anva16 TDn9a31 TDnva31 2e-014
Cn9anva17 TDn9a33 TDnva33 2e-014
Cn10an11a1 TDn10a1 TDn11a1 2e-014
Cn10an11a2 TDn10a3 TDn11a3 1e-014
Cn10an11a3 TDn10a5 TDn11a5 1e-014
Cn10an11a4 TDn10a7 TDn11a7 1e-014
Cn10an11a5 TDn10a9 TDn11a9 1e-014
Cn10an11a6 TDn10a11 TDn11a11 1e-014
Cn10an11a7 TDn10a13 TDn11a13 1e-014
Cn10an11a8 TDn10a15 TDn11a15 1e-014
Cn10an11a9 TDn10a17 TDn11a17 1e-014
Cn10an11a10 TDn10a19 TDn11a19 1e-014
Cn10an11a11 TDn10a21 TDn11a21 1e-014
Cn10an11a12 TDn10a23 TDn11a23 1e-014
Cn10an11a13 TDn10a25 TDn11a25 1e-014
Cn10an11a14 TDn10a27 TDn11a27 1e-014
Cn10an11a15 TDn10a29 TDn11a29 1e-014
Cn10an11a16 TDn10a31 TDn11a31 1e-014
Cn10an11a17 TDn10a33 TDn11a33 2e-014
Cn10an12a1 TDn10a1 TDn12a1 2e-014
Cn10an12a2 TDn10a3 TDn12a3 1e-014
Cn10an12a3 TDn10a5 TDn12a5 1e-014
Cn10an12a4 TDn10a7 TDn12a7 1e-014
Cn10an12a5 TDn10a9 TDn12a9 1e-014
Cn10an12a6 TDn10a11 TDn12a11 1e-014
Cn10an12a7 TDn10a13 TDn12a13 1e-014
Cn10an12a8 TDn10a15 TDn12a15 1e-014
Cn10an12a9 TDn10a17 TDn12a17 1e-014
Cn10an12a10 TDn10a19 TDn12a19 1e-014
Cn10an12a11 TDn10a21 TDn12a21 1e-014
Cn10an12a12 TDn10a23 TDn12a23 1e-014
Cn10an12a13 TDn10a25 TDn12a25 1e-014
Cn10an12a14 TDn10a27 TDn12a27 1e-014
Cn10an12a15 TDn10a29 TDn12a29 1e-014
Cn10an12a16 TDn10a31 TDn12a31 1e-014
Cn10an12a17 TDn10a33 TDn12a33 2e-014
Cn10anva1 TDn10a1 TDnva1 2e-014
Cn10anva2 TDn10a3 TDnva3 2e-014
Cn10anva3 TDn10a5 TDnva5 2e-014
Cn10anva4 TDn10a7 TDnva7 2e-014
Cn10anva5 TDn10a9 TDnva9 2e-014
Cn10anva6 TDn10a11 TDnva11 2e-014
Cn10anva7 TDn10a13 TDnva13 2e-014
Cn10anva8 TDn10a15 TDnva15 2e-014
Cn10anva9 TDn10a17 TDnva17 2e-014
Cn10anva10 TDn10a19 TDnva19 2e-014
Cn10anva11 TDn10a21 TDnva21 2e-014
Cn10anva12 TDn10a23 TDnva23 2e-014
Cn10anva13 TDn10a25 TDnva25 2e-014
Cn10anva14 TDn10a27 TDnva27 2e-014
Cn10anva15 TDn10a29 TDnva29 2e-014
Cn10anva16 TDn10a31 TDnva31 2e-014
Cn10anva17 TDn10a33 TDnva33 2e-014
Cn11an12a1 TDn11a1 TDn12a1 2e-014
Cn11an12a2 TDn11a3 TDn12a3 1e-014
Cn11an12a3 TDn11a5 TDn12a5 1e-014
Cn11an12a4 TDn11a7 TDn12a7 1e-014
Cn11an12a5 TDn11a9 TDn12a9 1e-014
Cn11an12a6 TDn11a11 TDn12a11 1e-014
Cn11an12a7 TDn11a13 TDn12a13 1e-014
Cn11an12a8 TDn11a15 TDn12a15 1e-014
Cn11an12a9 TDn11a17 TDn12a17 1e-014
Cn11an12a10 TDn11a19 TDn12a19 1e-014
Cn11an12a11 TDn11a21 TDn12a21 1e-014
Cn11an12a12 TDn11a23 TDn12a23 1e-014
Cn11an12a13 TDn11a25 TDn12a25 1e-014
Cn11an12a14 TDn11a27 TDn12a27 1e-014
Cn11an12a15 TDn11a29 TDn12a29 1e-014
Cn11an12a16 TDn11a31 TDn12a31 1e-014
Cn11an12a17 TDn11a33 TDn12a33 2e-014
Cn11anva1 TDn11a1 TDnva1 2e-014
Cn11anva2 TDn11a3 TDnva3 2e-014
Cn11anva3 TDn11a5 TDnva5 2e-014
Cn11anva4 TDn11a7 TDnva7 2e-014
Cn11anva5 TDn11a9 TDnva9 2e-014
Cn11anva6 TDn11a11 TDnva11 2e-014
Cn11anva7 TDn11a13 TDnva13 2e-014
Cn11anva8 TDn11a15 TDnva15 2e-014
Cn11anva9 TDn11a17 TDnva17 2e-014
Cn11anva10 TDn11a19 TDnva19 2e-014
Cn11anva11 TDn11a21 TDnva21 2e-014
Cn11anva12 TDn11a23 TDnva23 2e-014
Cn11anva13 TDn11a25 TDnva25 2e-014
Cn11anva14 TDn11a27 TDnva27 2e-014
Cn11anva15 TDn11a29 TDnva29 2e-014
Cn11anva16 TDn11a31 TDnva31 2e-014
Cn11anva17 TDn11a33 TDnva33 2e-014
Cn12anva1 TDn12a1 TDnva1 2e-014
Cn12anva2 TDn12a3 TDnva3 2e-014
Cn12anva3 TDn12a5 TDnva5 2e-014
Cn12anva4 TDn12a7 TDnva7 2e-014
Cn12anva5 TDn12a9 TDnva9 2e-014
Cn12anva6 TDn12a11 TDnva11 2e-014
Cn12anva7 TDn12a13 TDnva13 2e-014
Cn12anva8 TDn12a15 TDnva15 2e-014
Cn12anva9 TDn12a17 TDnva17 2e-014
Cn12anva10 TDn12a19 TDnva19 2e-014
Cn12anva11 TDn12a21 TDnva21 2e-014
Cn12anva12 TDn12a23 TDnva23 2e-014
Cn12anva13 TDn12a25 TDnva25 2e-014
Cn12anva14 TDn12a27 TDnva27 2e-014
Cn12anva15 TDn12a29 TDnva29 2e-014
Cn12anva16 TDn12a31 TDnva31 2e-014
Cn12anva17 TDn12a33 TDnva33 2e-014
.ENDS intercon

.AC		LIN		5000	0		30e+9
.PRINT  AC VR(TDN1a9) VI(TDN1a9)
.PROBE  V(TDN1a9)

.end
